* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP UP DOWN VCTRL CLK VDD FREERUN F6 VSS OUT LF CSVB EX
X0 a_23444_3994 a_22864_4398 VSS.t289 VSS.t288 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 VDD.t112 a_22948_2038 a_22864_2486 VDD.t111 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X2 a_23099_4907 a_23011_4951 VSS.t124 VSS.t123 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VSS.t301 a_23455_217 a_23407_261 VSS.t67 nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4 F6.t15 a_23423_n1258 VSS.t102 VSS.t101 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X5 OUT.t9 a_5840_7613.t1 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X6 a_22864_4398 a_22948_3950 a_22884_3994 VSS.t146 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7 VDD.t245 a_22388_2038.t2 a_22304_2486 VDD.t244 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X8 VCTRL.t19 FREERUN.t0 EX.t17 VSS.t153 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X9 a_n2908_12013 a_1220_12453 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X10 a_24891_4907 a_24803_4951 VSS.t155 VSS.t154 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X11 OUT.t10 a_5840_7613.t1 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X12 LF.t20 FREERUN.t1 VCTRL.t33 VDD.t157 pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.33u
X13 a_22539_3430 a_22451_3522 VDD.t22 VDD.t21 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 a_n558_2704.t1 a_11009_2840 a_14657_n1138 VSS.t40 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X15 VCTRL.t18 FREERUN.t2 EX.t16 VSS.t181 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X16 LF.t21 a_n17351_68.t2 VCTRL.t40 VSS.t196 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X17 a_22203_n358.t7 a_21855_n1258 VSS.t180 VSS.t179 nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
X18 VSS.t2 a_23455_1567 a_23407_1611 VSS.t1 nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X19 LF.t41 VSS.t152 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X20 a_21855_4398 CLK.t0 VSS.t112 VSS.t111 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X21 EX.t25 a_n17351_68.t3 VCTRL.t56 VDD.t212 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X22 EX.t26 a_n17351_68.t4 VCTRL.t57 VDD.t213 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X23 VCTRL.t58 a_n17351_68.t5 EX.t27 VDD.t214 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X24 a_25265_7733 a_24755_6933 OUT.t7 VDD.t260 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X25 a_22203_n358.t6 a_21855_n1258 VSS.t178 VSS.t177 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X26 VSS.t100 a_23423_n1258 F6.t14 VSS.t99 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X27 VCTRL.t71 a_n17351_68.t6 EX.t32 VDD.t241 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X28 VSS.t260 a_n4208_n141.t3 a_n671_n1138 VSS.t259 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X29 VDD.t228 a_n8471_219.t5 a_3149_2840 VDD.t227 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X30 a_21755_1082 a_24383_1567 VSS.t49 VSS.t48 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X31 EX.t33 a_n17351_68.t7 VCTRL.t72 VDD.t242 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X32 VDD.t283 a_23620_8319.t3 a_23691_7733 VDD.t282 pfet_03v3 ad=1.3p pd=5.3u as=0.52p ps=2.52u w=2u l=0.33u
X33 VCTRL.t32 FREERUN.t3 LF.t19 VDD.t158 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X34 VSS.t68 a_23455_n345 a_23407_n301 VSS.t67 nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X35 VSS.t131 a_n8537_n1530.t4 a_n8659_n1230 VSS.t130 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X36 a_22987_3430 a_22899_3522 VDD.t97 VDD.t96 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X37 a_25675_477 a_25587_574 VSS.t211 VSS.t210 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X38 VDD.t225 a_22203_n358.t8 a_22115_253.t0 VDD.t224 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X39 a_7177_2840 a_3345_2840 a_6981_2840 VDD.t41 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X40 VDD.t13 a_23508_2038 a_22948_2038 VDD.t12 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X41 a_27014_14933 a_24866_11400 VSS.t45 ppolyf_u r_width=0.8u r_length=22u
X42 LF.t42 VSS.t209 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X43 VCTRL.t73 a_n17351_68.t8 EX.t34 VDD.t243 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X44 VDD.t156 a_21855_n1258 a_22203_n358.t3 VDD.t155 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X45 a_22948_3950 a_23508_2038 a_23444_3994 VSS.t10 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X46 OUT.t11 a_5840_7613.t1 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X47 a_26795_6933 a_n8537_93.t3 a_25265_6933 VSS.t267 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X48 EX.t38 a_n17351_68.t9 VCTRL.t77 VDD.t315 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X49 a_1220_13333 a_5840_13333 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X50 LF.t40 a_n17351_68.t10 VCTRL.t78 VSS.t300 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X51 VDD.t191 CSVB.t14 CSVB.t15 VDD.t190 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X52 a_24383_217 a_24090_629 VDD.t133 VDD.t132 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X53 VCTRL.t79 a_n17351_68.t11 EX.t39 VDD.t316 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X54 a_1712_14653 OUT.t3 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X55 VSS.t217 a_16431_6193 VSS.t13 ppolyf_u r_width=0.8u r_length=0.13m
X56 a_23407_1611 a_22527_1197 a_23083_1611 VSS.t20 nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X57 a_21643_3430 a_21555_3522 VDD.t262 VDD.t261 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X58 a_n8471_219.t4 a_n8537_93.t4 a_n8659_n1230 VSS.t268 nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.33u
X59 a_26049_6873 DOWN.t2 VDD.t309 VDD.t308 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X60 a_22864_4398 a_22304_4398 VDD.t94 VDD.t93 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X61 a_21506_13215.t9 CSVB.t18 VDD.t198 VDD.t197 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X62 a_23083_1611 a_22963_1518 a_22915_1611 VSS.t242 nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X63 VCTRL.t31 FREERUN.t4 LF.t18 VDD.t141 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X64 a_n2908_11133 a_1220_11573 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X65 a_22304_4398 a_21855_4398 VDD.t3 VDD.t2 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X66 EX.t20 a_n17351_68.t12 VCTRL.t41 VDD.t176 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X67 VCTRL.t42 a_n17351_68.t13 LF.t22 VSS.t204 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X68 VSS.t110 UP.t2 a_24755_6933 VSS.t109 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X69 F6.t7 a_23423_n1258 VDD.t81 VDD.t80 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X70 VDD.t230 a_n8471_219.t6 a_18477_2840 VDD.t229 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X71 VDD.t277 a_22864_2486 a_22388_2038.t1 VDD.t276 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X72 VDD.t79 a_23423_n1258 F6.t6 VDD.t78 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X73 VCTRL.t43 a_n17351_68.t14 EX.t21 VDD.t177 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X74 a_23083_261 a_22963_217 a_22915_261 VSS.t35 nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X75 VSS.t218 a_25675_n394 a_25587_n302 VSS.t210 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X76 a_22959_n669 a_22527_n715 VDD.t205 VDD.t204 pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X77 VSS.t98 a_23423_n1258 F6.t13 VSS.t97 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X78 VDD.t207 CSVB.t19 a_21506_13215.t8 VDD.t206 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X79 a_23407_n301 a_22527_n715 a_23083_n301 VSS.t74 nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X80 a_21855_1126 a_21755_1082 VSS.t64 VSS.t62 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X81 a_21855_n1258 a_n558_2704.t2 VSS.t172 VSS.t171 nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X82 EX.t35 a_n17351_68.t15 VCTRL.t74 VDD.t269 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X83 a_22959_1243 a_22527_1197 VDD.t20 VDD.t19 pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X84 VSS.t133 a_n8537_n1530.t5 a_21891_6933 VSS.t132 nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.33u
X85 LF.t43 VSS.t106 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X86 EX.t36 a_n17351_68.t16 VCTRL.t75 VDD.t270 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X87 a_25265_7733 a_22941_7733.t3 a_25095_7733 VDD.t136 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X88 a_23083_n301 a_21855_1126 a_22915_n301 VSS.t35 nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X89 OUT.t12 a_5840_7613.t1 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X90 VCTRL.t76 a_n17351_68.t17 EX.t37 VDD.t271 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X91 VSS.t246 a_n8537_n1530.t6 a_n8659_n1230 VSS.t245 nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.33u
X92 LF.t38 a_n17351_68.t18 VCTRL.t68 VSS.t240 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X93 LF.t17 FREERUN.t5 VCTRL.t22 VDD.t142 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X94 a_22941_7733.t2 a_n8537_93.t5 a_22955_6933 VSS.t243 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X95 a_24383_n345 a_24090_n669 VDD.t170 VDD.t169 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X96 a_23427_629 a_22115_253.t2 a_23083_261 VDD.t86 pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X97 a_21755_1082 a_24383_1567 VDD.t34 VDD.t33 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X98 a_22527_1197 a_22115_1610.t2 VSS.t32 VSS.t31 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X99 VDD.t226 a_22203_n358.t9 a_22115_1610.t0 VDD.t224 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X100 a_21855_n1258 a_n558_2704.t3 VDD.t188 VDD.t187 pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X101 a_21506_13215.t7 CSVB.t20 VDD.t209 VDD.t208 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X102 VCTRL.t17 FREERUN.t6 EX.t1 VSS.t167 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X103 F6.t12 a_23423_n1258 VSS.t96 VSS.t95 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X104 a_22527_574 a_22115_253.t3 VDD.t87 VDD.t82 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X105 a_23083_n301 a_21855_1126 a_22959_n669 VDD.t27 pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X106 VSS.t61 a_22091_3430 a_22003_3522 VSS.t60 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X107 a_26115_6933 a_26049_6873 a_25265_6933 VSS.t24 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X108 a_23407_261 a_22527_574 a_23083_261 VSS.t74 nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X109 a_23083_1611 a_22963_1518 a_22959_1243 VDD.t246 pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X110 a_22915_1611 a_22115_1610.t3 VSS.t34 VSS.t33 nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X111 a_22948_3950 a_22864_4398 VDD.t297 VDD.t296 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X112 VCTRL.t21 FREERUN.t7 LF.t16 VDD.t162 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X113 a_22203_n358.t2 a_21855_n1258 VDD.t154 VDD.t153 pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X114 a_23435_3430 a_23347_3522 VDD.t46 VDD.t45 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X115 EX.t31 a_n17351_68.t19 VCTRL.t69 VDD.t240 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X116 VCTRL.t70 a_n17351_68.t20 LF.t39 VSS.t241 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X117 VDD.t275 a_22864_2486 a_23508_2038 VDD.t274 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X118 a_24207_4398 a_22304_4398 VSS.t119 VSS.t118 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X119 a_23455_217 a_23083_261 VSS.t6 VSS.t5 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X120 VDD.t266 a_n8471_219.t0 a_n8471_219.t1 VDD.t265 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X121 a_25265_7733 UP.t3 a_26115_6933 VDD.t14 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X122 a_23423_n1258 a_22203_n358.t10 VSS.t230 VSS.t229 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X123 EX.t0 FREERUN.t8 VCTRL.t16 VSS.t188 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X124 a_22203_n358.t1 a_21855_n1258 VDD.t152 VDD.t151 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X125 VDD.t192 a_25675_477 a_25587_574 VDD.t134 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X126 F6.t5 a_23423_n1258 VDD.t77 VDD.t76 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X127 a_22915_n301 a_22115_n302.t2 VSS.t252 VSS.t113 nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X128 a_23423_n1258 a_22203_n358.t11 VSS.t232 VSS.t231 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X129 VDD.t317 a_23455_217 a_23427_629 VDD.t0 pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X130 LF.t44 VSS.t107 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X131 a_23691_7733 a_23620_8319.t4 VDD.t36 VDD.t35 pfet_03v3 ad=0.52p pd=2.52u as=1.3p ps=5.3u w=2u l=0.33u
X132 a_n2908_7613 VSS.t44 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X133 a_22388_3950.t1 a_23508_2038 VDD.t11 VDD.t10 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X134 LF.t15 FREERUN.t9 VCTRL.t20 VDD.t163 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X135 VSS.t248 a_n8537_n1530.t7 a_22955_6933 VSS.t247 nfet_03v3 ad=0.4p pd=1.8u as=0.26p ps=1.52u w=1u l=0.33u
X136 a_n2908_10253 a_1220_10693 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X137 a_23883_3430 a_23795_3522 VDD.t85 VDD.t84 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X138 a_24655_4398 a_24207_4398 VSS.t57 VSS.t56 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X139 a_n2908_9373 a_1220_8933 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X140 VDD.t26 a_21755_4907 a_21667_4951 VDD.t25 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X141 a_21855_4398 CLK.t1 VDD.t140 VDD.t139 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X142 a_22388_3950.t1 a_24655_4398 VDD.t256 VDD.t255 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X143 VCTRL.t15 FREERUN.t10 EX.t13 VSS.t182 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X144 a_21755_477 a_21667_574 VSS.t148 VSS.t147 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X145 a_11009_2840 a_7177_2840 a_10813_2840 VDD.t249 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X146 VDD.t232 a_n8471_219.t7 a_n683_2840 VDD.t231 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X147 UP.t0 a_22388_3950.t2 VSS.t166 VSS.t165 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X148 EX.t28 a_n17351_68.t21 VCTRL.t59 VDD.t216 pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.33u
X149 LF.t32 a_n17351_68.t22 VCTRL.t60 VSS.t225 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X150 a_26115_6933 a_26049_6873 a_25265_6933 VSS.t23 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X151 a_25150_3994 a_24655_4398 VSS.t256 VSS.t255 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X152 a_22304_4398 a_22388_3950.t3 a_22324_3994 VSS.t279 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X153 VSS.t176 a_21855_n1258 a_22203_n358.t5 VSS.t175 nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X154 VCTRL.t14 FREERUN.t11 EX.t12 VSS.t183 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X155 VCTRL.t25 FREERUN.t12 LF.t14 VDD.t159 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X156 a_21506_13215.t6 CSVB.t21 VDD.t211 VDD.t210 pfet_03v3 ad=1.456p pd=6.12u as=3.64p ps=12.5u w=5.6u l=0.56u
X157 VSS.t234 a_22203_n358.t12 a_22115_1610.t1 VSS.t233 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X158 a_22963_217 a_24383_n345 VDD.t56 VDD.t55 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X159 a_25265_7733 UP.t4 a_26115_6933 VDD.t15 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X160 a_22388_2038.t0 a_23508_2038 a_25334_2082 VSS.t9 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X161 a_23620_8319.t2 a_n8537_93.t6 a_23691_6933 VSS.t244 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X162 VDD.t144 CSVB.t22 a_21506_13215.t5 VDD.t143 pfet_03v3 ad=3.64p pd=12.5u as=1.456p ps=6.12u w=5.6u l=0.56u
X163 a_1712_7613 a_5840_7613.t0 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X164 VDD.t281 a_22941_7733.t0 a_22941_7733.t1 VDD.t280 pfet_03v3 ad=1.072p pd=5.3u as=1.072p ps=5.3u w=0.8u l=0.33u
X165 VDD.t264 a_24383_217 a_24375_629 VDD.t31 pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X166 VCTRL.t61 a_n17351_68.t23 LF.t33 VSS.t226 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X167 VDD.t200 a_n558_2704.t4 a_21855_n1258 VDD.t199 pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X168 a_1712_9373 a_5840_8933 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X169 a_23691_7733 a_22941_7733.t4 a_23620_8319.t1 VDD.t137 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X170 a_21891_6933 a_n8537_n1530.t8 VSS.t84 VSS.t83 nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.33u
X171 a_1712_11133 a_5840_11573 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X172 a_n2908_14213 a_1220_14653 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X173 a_24755_6933 UP.t5 VDD.t254 VDD.t253 pfet_03v3 ad=0.52p pd=2.52u as=1.3p ps=5.3u w=2u l=0.33u
X174 a_22915_261 a_22115_253.t4 VSS.t114 VSS.t113 nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X175 a_24090_629 a_22115_253.t5 a_23455_217 VDD.t88 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X176 OUT.t13 a_5840_7613.t1 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X177 LF.t29 a_n17351_68.t24 VCTRL.t53 VSS.t222 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X178 VDD.t146 CSVB.t23 a_21506_13215.t4 VDD.t145 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X179 VCTRL.t24 FREERUN.t13 LF.t13 VDD.t193 pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.33u
X180 LF.t12 FREERUN.t14 VCTRL.t23 VDD.t194 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X181 VDD.t30 a_23547_4907 a_23459_4951 VDD.t29 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X182 VSS.t278 a_n8537_93.t1 a_n8537_93.t2 VSS.t277 nfet_03v3 ad=0.496p pd=3.22u as=0.496p ps=3.22u w=0.4u l=0.33u
X183 VSS.t237 a_22203_n358.t13 a_23423_n1258 VSS.t236 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X184 a_27814_14933 a_27414_10401 VSS.t104 ppolyf_u r_width=0.8u r_length=22u
X185 a_25104_3522 a_22304_4398 a_24900_3522 VSS.t117 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X186 a_3345_2840 a_n487_2840 a_3149_2840 VDD.t95 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X187 OUT.t14 a_5840_7613.t1 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X188 a_25334_3994 a_22864_4398 a_25150_3994 VSS.t287 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X189 a_22884_2082 a_22304_2486 VSS.t80 VSS.t79 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X190 a_22527_574 a_22115_253.t6 VSS.t302 VSS.t290 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X191 VDD.t38 a_23620_8319.t5 a_26795_7733 VDD.t37 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X192 a_n2908_8493 a_1220_8053 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X193 a_25265_6933 DOWN.t3 OUT.t1 VSS.t140 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X194 LF.t45 VSS.t152 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X195 a_22324_2082 a_21855_2486 VSS.t285 VSS.t284 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X196 a_7177_2840 a_3345_2840 a_6993_n1138 VSS.t58 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X197 a_n487_2840 a_n558_2704.t5 a_n671_n1138 VSS.t197 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X198 OUT.t15 a_5840_7613.t1 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X199 CSVB.t13 CSVB.t12 VDD.t121 VDD.t120 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X200 a_24335_261 a_22115_253.t7 a_24090_629 VSS.t164 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X201 a_23455_n345 a_23083_n301 VDD.t131 VDD.t130 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X202 VDD.t182 a_22203_4907 a_22115_4951 VDD.t181 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X203 OUT.t6 a_24755_6933 a_25265_7733 VDD.t259 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X204 a_22527_n715 a_22115_n302.t3 VDD.t252 VDD.t251 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X205 VDD.t165 a_23995_4907 a_23907_4951 VDD.t164 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X206 a_23455_1567 a_23083_1611 VDD.t250 VDD.t4 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X207 a_n4208_n141.t2 a_n8471_219.t8 VDD.t219 VDD.t218 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X208 LF.t11 FREERUN.t15 VCTRL.t39 VDD.t195 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X209 F6.t4 a_23423_n1258 VDD.t75 VDD.t74 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X210 VSS.t94 a_23423_n1258 F6.t11 VSS.t93 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X211 a_23455_217 a_23083_261 VDD.t5 VDD.t4 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X212 VDD.t268 a_21755_477 a_21667_574 VDD.t267 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X213 a_22955_6933 a_n8537_n1530.t9 VSS.t86 VSS.t85 nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.33u
X214 LF.t46 VSS.t209 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X215 a_1712_8493 a_5840_8053 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X216 a_24207_4398 a_22304_4398 VDD.t92 VDD.t91 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X217 VSS.t16 a_25675_1518 a_25587_1610 VSS.t15 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X218 a_21855_2486 a_21755_1082 VSS.t63 VSS.t62 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X219 VDD.t99 a_22651_4907 a_22563_4951 VDD.t98 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X220 a_23444_2082 a_22864_2486 VSS.t266 VSS.t265 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X221 VDD.t105 a_25339_4907 a_25251_4951 VDD.t104 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X222 a_18673_2840 a_n558_2704.t6 a_18477_2840 VDD.t215 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X223 a_1712_10253 a_5840_10693 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X224 a_24383_217 a_24090_629 VSS.t151 VSS.t150 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X225 a_n2908_13333 a_1220_13773 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X226 VCTRL.t54 a_n17351_68.t25 LF.t30 VSS.t223 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X227 a_25265_6933 DOWN.t4 OUT.t2 VSS.t141 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X228 VDD.t150 a_21855_n1258 a_22203_n358.t0 VDD.t149 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X229 VDD.t52 a_23455_n345 a_23427_n669 VDD.t51 pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X230 EX.t3 FREERUN.t16 VCTRL.t13 VSS.t184 nfet_03v3 ad=0.26p pd=1.52u as=0.65p ps=3.3u w=1u l=0.33u
X231 a_21855_1126 a_21755_1082 VDD.t50 VDD.t49 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X232 a_22864_2486 a_22948_2038 a_22884_2082 VSS.t127 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X233 VSS.t135 a_n8537_n1530.t10 a_23691_6933 VSS.t134 nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.33u
X234 VDD.t1 a_23455_1567 a_23427_1243 VDD.t0 pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X235 a_23508_2038 a_22304_2486 VDD.t63 VDD.t62 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X236 a_n8471_219.t3 VCTRL.t80 a_n9701_6193 VSS.t274 nfet_03v3 ad=0.488p pd=2.82u as=0.488p ps=2.82u w=0.8u l=0.33u
X237 EX.t2 FREERUN.t17 VCTRL.t12 VSS.t185 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X238 a_18673_2840 a_n558_2704.t7 a_18489_n1138 VSS.t216 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X239 a_24655_4398 a_24207_4398 VDD.t40 VDD.t39 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X240 VDD.t234 a_22203_n358.t14 a_23423_n1258 VDD.t233 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X241 LF.t10 FREERUN.t18 VCTRL.t38 VDD.t160 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
D0 VSS.t129 VSS.t128 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X242 a_n2908_12013 a_1220_11573 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X243 a_24383_1567 a_24090_1243 VSS.t299 VSS.t298 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X244 UP.t1 a_22388_3950.t4 VDD.t289 VDD.t288 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X245 EX.t19 FREERUN.t19 VCTRL.t11 VSS.t168 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X246 a_23508_2038 a_22864_4398 a_25104_3522 VSS.t286 nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X247 a_25095_7733 a_23620_8319.t6 VDD.t301 VDD.t300 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X248 a_23455_1567 a_23083_1611 VSS.t251 VSS.t250 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X249 a_22091_3430 a_22003_3522 VDD.t17 VDD.t16 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X250 a_24866_11400 a_21506_13215.t10 CSVB.t16 VSS.t38 nfet_03v3 ad=3.416p pd=12.42u as=1.456p ps=6.12u w=5.6u l=0.56u
X251 VCTRL.t10 FREERUN.t20 EX.t18 VSS.t169 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X252 a_26049_6873 DOWN.t5 VSS.t126 VSS.t125 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X253 a_22959_629 a_22527_574 VDD.t57 VDD.t19 pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X254 a_22864_2486 a_22304_2486 VDD.t61 VDD.t60 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X255 VSS.t262 a_n4208_n141.t4 a_18489_n1138 VSS.t261 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X256 a_24383_n345 a_24090_n669 VSS.t198 VSS.t150 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X257 VCTRL.t55 a_n17351_68.t26 LF.t31 VSS.t224 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X258 VDD.t73 a_23423_n1258 F6.t3 VDD.t72 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X259 a_22304_2486 a_21855_2486 VDD.t291 VDD.t290 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X260 VDD.t24 a_24443_4907 a_24355_4951 VDD.t23 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X261 VCTRL.t9 FREERUN.t21 EX.t11 VSS.t170 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X262 a_1712_14653 a_5840_14213 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X263 VDD.t103 DOWN.t6 a_26049_6873 VDD.t102 pfet_03v3 ad=1.3p pd=5.3u as=0.52p ps=2.52u w=2u l=0.33u
X264 a_22948_2038 a_23508_2038 a_23444_2082 VSS.t8 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X265 VDD.t295 a_22864_4398 a_23508_2038 VDD.t294 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X266 a_23455_n345 a_23083_n301 VSS.t149 VSS.t5 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X267 OUT.t16 a_5840_7613.t1 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X268 a_24383_1567 a_24090_1243 VDD.t314 VDD.t132 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X269 VCTRL.t8 FREERUN.t22 EX.t10 VSS.t296 nfet_03v3 ad=0.65p pd=3.3u as=0.26p ps=1.52u w=1u l=0.33u
X270 a_25265_6933 a_n8537_93.t7 a_25095_6933 VSS.t303 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X271 LF.t9 FREERUN.t23 VCTRL.t37 VDD.t312 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X272 a_n2908_9373 a_1220_9813 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X273 VDD.t319 a_23099_4907 a_23011_4951 VDD.t318 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X274 VDD.t117 a_21755_n830 a_21667_n786 VDD.t116 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X275 a_n487_2840 a_n558_2704.t8 a_n683_2840 VDD.t189 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X276 OUT.t5 a_24755_6933 a_25265_7733 VDD.t258 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X277 VDD.t248 a_24891_4907 a_24803_4951 VDD.t247 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X278 CSVB.t11 CSVB.t10 VDD.t119 VDD.t118 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X279 LF.t23 a_n17351_68.t27 VCTRL.t47 VSS.t206 nfet_03v3 ad=0.26p pd=1.52u as=0.65p ps=3.3u w=1u l=0.33u
X280 VDD.t54 a_24383_n345 a_24375_n669 VDD.t53 pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X281 VCTRL.t28 FREERUN.t24 LF.t8 VDD.t313 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X282 a_22955_6933 a_n8537_93.t8 a_22941_7733.t2 VSS.t304 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X283 VDD.t32 a_24383_1567 a_24375_1243 VDD.t31 pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X284 a_24375_629 a_22527_574 a_24090_629 VDD.t18 pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X285 a_22948_2038 a_22864_2486 VDD.t273 VDD.t272 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X286 a_n2908_11133 a_1220_10693 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X287 a_24207_2486 a_22304_2486 VSS.t78 VSS.t77 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X288 LF.t47 VSS.t108 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X289 VDD.t311 CSVB.t8 CSVB.t9 VDD.t310 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X290 a_25265_6933 a_26049_6873 a_26115_6933 VSS.t22 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X291 a_22963_1518 a_24383_217 VSS.t258 VSS.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X292 a_1712_9373 a_5840_9813 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X293 VDD.t127 a_22948_3950 a_22864_4398 VDD.t126 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X294 LF.t7 FREERUN.t25 VCTRL.t27 VDD.t201 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X295 VSS.t39 a_24866_11400 a_21506_13215.t1 VSS.t38 nfet_03v3 ad=3.416p pd=12.42u as=1.456p ps=6.12u w=5.6u l=0.56u
X296 a_n8659_n1230 a_n8537_n1530.t11 VSS.t137 VSS.t136 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X297 VCTRL.t48 a_n17351_68.t28 LF.t24 VSS.t207 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X298 VDD.t287 a_22388_3950.t5 a_22304_4398 VDD.t286 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X299 a_24335_1611 a_22115_1610.t4 a_24090_1243 VSS.t103 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X300 a_23691_6933 a_n8537_n1530.t12 VSS.t28 VSS.t27 nfet_03v3 ad=0.26p pd=1.52u as=0.4p ps=1.8u w=1u l=0.33u
X301 a_22388_2038.t1 a_23508_2038 VDD.t9 VDD.t8 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X302 EX.t9 FREERUN.t26 VCTRL.t7 VSS.t221 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X303 CSVB.t7 CSVB.t6 VDD.t125 VDD.t124 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X304 a_1712_13773 a_5840_13333 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X305 a_24655_2486 a_24207_2486 VSS.t143 VSS.t142 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X306 a_24090_1243 a_22527_1197 a_23455_1567 VSS.t19 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X307 a_21855_2486 a_21755_1082 VDD.t48 VDD.t47 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X308 a_22388_2038.t1 a_24655_2486 VDD.t65 VDD.t64 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X309 VDD.t148 CSVB.t24 a_21506_13215.t3 VDD.t147 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X310 F6.t10 a_23423_n1258 VSS.t92 VSS.t91 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X311 VCTRL.t26 FREERUN.t27 LF.t6 VDD.t202 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X312 DOWN.t1 a_22388_2038.t3 VSS.t139 VSS.t138 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X313 a_22963_1518 a_24383_217 VDD.t263 VDD.t33 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X314 VSS.t190 a_n4208_n141.t5 a_14657_n1138 VSS.t189 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X315 a_24335_n301 a_22115_n302.t4 a_24090_n669 VSS.t164 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X316 a_22527_1197 a_22115_1610.t5 VDD.t83 VDD.t82 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X317 a_n2908_8493 a_1220_8933 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X318 VCTRL.t6 FREERUN.t28 EX.t8 VSS.t186 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X319 a_1220_12453 a_5840_11573 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X320 VDD.t221 a_n8471_219.t9 a_14645_2840 VDD.t220 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X321 a_23427_n669 a_22115_n302.t5 a_23083_n301 VDD.t138 pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X322 VCTRL.t49 a_n17351_68.t29 LF.t25 VSS.t208 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X323 a_25265_6933 a_26049_6873 a_26115_6933 VSS.t21 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X324 a_23083_261 a_22963_217 a_22959_629 VDD.t246 pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X325 a_24090_n669 a_22527_n715 a_23455_n345 VSS.t73 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X326 a_23427_1243 a_22115_1610.t6 a_23083_1611 VDD.t86 pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X327 VDD.t7 a_23508_2038 a_22948_3950 VDD.t6 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X328 a_23508_2038 a_22304_4398 VDD.t90 VDD.t89 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X329 a_26795_7733 a_22941_7733.t5 a_25265_7733 VDD.t284 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X330 a_23691_6933 a_n8537_93.t9 a_23620_8319.t0 VSS.t156 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X331 a_n2908_10253 a_1220_9813 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X332 a_21755_4907 a_21667_4951 VSS.t145 VSS.t144 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X333 OUT.t17 a_5840_7613.t1 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X334 a_25150_2082 a_24655_2486 VSS.t82 VSS.t81 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X335 a_22304_2486 a_22388_2038.t4 a_22324_2082 VSS.t235 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X336 EX.t5 FREERUN.t29 VCTRL.t5 VSS.t187 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X337 LF.t5 FREERUN.t30 VCTRL.t36 VDD.t161 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X338 VDD.t236 a_22203_n358.t15 a_23423_n1258 VDD.t235 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X339 OUT.t18 a_5840_7613.t1 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X340 VSS.t192 a_n4208_n141.t6 a_3161_n1138 VSS.t191 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X341 a_27014_14933 a_27414_10401 VSS.t59 ppolyf_u r_width=0.8u r_length=22u
X342 LF.t26 a_n17351_68.t30 VCTRL.t50 VSS.t213 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X343 a_24755_6933 UP.t6 VSS.t254 VSS.t253 nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.33u
X344 a_1712_8493 a_5840_8933 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X345 VSS.t12 a_22539_3430 a_22451_3522 VSS.t11 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X346 EX.t4 FREERUN.t31 VCTRL.t4 VSS.t294 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X347 a_25675_1518 a_25587_1610 VDD.t135 VDD.t134 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X348 CSVB.t5 CSVB.t4 VDD.t123 VDD.t122 pfet_03v3 ad=1.456p pd=6.12u as=3.64p ps=12.5u w=5.6u l=0.56u
X349 a_21891_6933 a_n8537_93.t10 a_n8537_n1530.t0 VSS.t157 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X350 VDD.t43 UP.t7 a_24755_6933 VDD.t42 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X351 CSVB.t17 a_21506_13215.t11 a_24866_11400 VSS.t36 nfet_03v3 ad=1.456p pd=6.12u as=3.416p ps=12.42u w=5.6u l=0.56u
X352 VDD.t293 a_22864_4398 a_22388_3950.t1 VDD.t292 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X353 VDD.t129 CSVB.t2 CSVB.t3 VDD.t128 pfet_03v3 ad=3.64p pd=12.5u as=1.456p ps=6.12u w=5.6u l=0.56u
X354 VCTRL.t51 a_n17351_68.t31 LF.t27 VSS.t214 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X355 VSS.t30 a_n8537_n1530.t13 a_26795_6933 VSS.t29 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X356 VCTRL.t35 FREERUN.t32 LF.t4 VDD.t299 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X357 VSS.t200 a_22203_n358.t16 a_22115_253.t1 VSS.t199 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X358 a_n4208_n141.t1 a_n4208_n141.t0 VSS.t122 VSS.t121 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X359 VCTRL.t3 FREERUN.t33 EX.t7 VSS.t295 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X360 VSS.t66 a_22987_3430 a_22899_3522 VSS.t65 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X361 a_22963_217 a_24383_n345 VSS.t72 VSS.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X362 a_n8471_219.t2 a_n8537_93.t11 a_n8659_n1230 VSS.t25 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X363 a_24090_629 a_22527_574 a_23455_217 VSS.t73 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X364 VDD.t223 a_n8471_219.t10 a_6981_2840 VDD.t222 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X365 OUT.t8 DOWN.t7 a_25265_6933 VSS.t269 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X366 VDD.t71 a_23423_n1258 F6.t2 VDD.t70 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X367 VSS.t90 a_23423_n1258 F6.t9 VSS.t89 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X368 a_1712_11133 a_5840_10693 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X369 LF.t3 FREERUN.t34 VCTRL.t34 VDD.t166 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X370 a_n2908_14213 a_1220_13773 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
D1 VSS.t305 VDD.t113 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X371 a_n17351_68.t0 FREERUN.t35 VDD.t168 VDD.t167 pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.28u
X372 LF.t28 a_n17351_68.t32 VCTRL.t52 VSS.t215 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X373 VDD.t186 CSVB.t0 CSVB.t1 VDD.t185 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X374 VDD.t303 CSVB.t25 a_n8537_n1530.t2 VDD.t302 pfet_03v3 ad=1.456p pd=5.78u as=0.5824p ps=2.76u w=2.24u l=0.56u
X375 a_23547_4907 a_23459_4951 VSS.t55 VSS.t54 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X376 a_25334_2082 a_22864_2486 a_25150_2082 VSS.t264 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X377 a_26115_6933 UP.t8 a_25265_7733 VDD.t44 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X378 VSS.t47 a_24383_1567 a_24335_1611 VSS.t46 nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X379 EX.t6 FREERUN.t36 VCTRL.t2 VSS.t195 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X380 VSS.t159 a_21643_3430 a_21555_3522 VSS.t158 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X381 a_11009_2840 a_7177_2840 a_10825_n1138 VSS.t249 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X382 a_24207_2486 a_22304_2486 VDD.t59 VDD.t58 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X383 LF.t48 VSS.t106 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X384 a_24706_3522 a_22304_2486 VSS.t76 VSS.t75 nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X385 VSS.t194 a_n4208_n141.t7 a_6993_n1138 VSS.t193 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X386 a_23423_n1258 a_22203_n358.t17 VDD.t172 VDD.t171 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X387 VCTRL.t65 a_n17351_68.t33 LF.t36 VSS.t238 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X388 a_n2908_7613 a_1220_8053 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X389 VSS.t70 a_24383_n345 a_24335_n301 VSS.t69 nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X390 a_22203_4907 a_22115_4951 VSS.t283 VSS.t282 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X391 a_25675_n394 a_25587_n302 VDD.t101 VDD.t100 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X392 OUT.t19 VSS.t43 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X393 a_23423_n1258 a_22203_n358.t18 VDD.t174 VDD.t173 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X394 a_23995_4907 a_23907_4951 VSS.t281 VSS.t280 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X395 a_24375_n669 a_22527_n715 a_24090_n669 VDD.t203 pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X396 a_22388_3950.t0 a_23508_2038 a_25334_3994 VSS.t7 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X397 a_24375_1243 a_22527_1197 a_24090_1243 VDD.t18 pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X398 a_n8537_n1530.t3 CSVB.t26 VDD.t305 VDD.t304 pfet_03v3 ad=0.5824p pd=2.76u as=0.5824p ps=2.76u w=2.24u l=0.56u
X399 a_21506_13215.t0 a_24866_11400 VSS.t37 VSS.t36 nfet_03v3 ad=1.456p pd=6.12u as=3.416p ps=12.42u w=5.6u l=0.56u
X400 a_24655_2486 a_24207_2486 VDD.t115 VDD.t114 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X401 a_21755_n830 a_21667_n786 VSS.t297 VSS.t147 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X402 a_n8659_n1230 a_n8537_n1530.t14 VSS.t161 VSS.t160 nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.33u
X403 a_n8659_n1230 a_n8537_93.t12 a_n8471_219.t2 VSS.t26 nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.33u
X404 a_24900_3522 a_22864_2486 a_24706_3522 VSS.t263 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X405 F6.t1 a_23423_n1258 VDD.t69 VDD.t68 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X406 DOWN.t0 a_22388_2038.t5 VDD.t279 VDD.t278 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X407 a_26115_6933 UP.t9 a_25265_7733 VDD.t106 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X408 VDD.t67 a_23423_n1258 F6.t0 VDD.t66 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X409 OUT.t20 a_5840_7613.t1 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X410 a_27814_14933 VSS.t53 VSS.t52 ppolyf_u r_width=0.8u r_length=22u
X411 VCTRL.t66 a_n17351_68.t34 EX.t30 VDD.t239 pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.33u
X412 a_22651_4907 a_22563_4951 VSS.t273 VSS.t272 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X413 a_25095_6933 a_n8537_n1530.t15 VSS.t163 VSS.t162 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X414 a_22527_n715 a_22115_n302.t6 VSS.t291 VSS.t290 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X415 a_1712_7613 a_5840_8053 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X416 VCTRL.t30 FREERUN.t37 LF.t2 VDD.t175 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X417 a_25339_4907 a_25251_4951 VSS.t42 VSS.t41 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X418 VSS.t220 a_n4208_n141.t8 a_10825_n1138 VSS.t219 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X419 VCTRL.t67 a_n17351_68.t35 LF.t37 VSS.t239 nfet_03v3 ad=0.65p pd=3.3u as=0.26p ps=1.52u w=1u l=0.33u
X420 LF.t34 a_n17351_68.t36 VCTRL.t62 VSS.t227 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X421 a_3345_2840 a_n487_2840 a_3161_n1138 VSS.t120 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X422 a_1712_10253 a_5840_9813 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X423 a_n8537_93.t0 CSVB.t27 VDD.t307 VDD.t306 pfet_03v3 ad=0.5824p pd=2.76u as=1.456p ps=5.78u w=2.24u l=0.56u
X424 a_23620_8319.t1 a_22941_7733.t6 a_23691_7733 VDD.t285 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X425 VDD.t184 a_22203_n358.t19 a_22115_n302.t0 VDD.t183 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X426 a_n2908_13333 a_1220_13333 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X427 VSS.t18 a_23435_3430 a_23347_3522 VSS.t17 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X428 LF.t49 VSS.t107 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X429 a_24090_n669 a_22115_n302.t7 a_23455_n345 VDD.t298 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X430 VSS.t174 a_21855_n1258 a_22203_n358.t4 VSS.t173 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X431 F6.t8 a_23423_n1258 VSS.t88 VSS.t87 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X432 VSS.t271 DOWN.t8 a_26049_6873 VSS.t270 nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.33u
X433 LF.t0 a_1220_14653 VSS.t14 ppolyf_u_1k r_width=1u r_length=20u
X434 VDD.t108 CSVB.t28 a_n8537_93.t0 VDD.t107 pfet_03v3 ad=0.5824p pd=2.76u as=0.5824p ps=2.76u w=2.24u l=0.56u
X435 a_22884_3994 a_22304_4398 VSS.t116 VSS.t115 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X436 LF.t50 VSS.t108 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X437 a_24090_1243 a_22115_1610.t7 a_23455_1567 VDD.t88 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X438 a_21506_13215.t2 CSVB.t29 VDD.t110 VDD.t109 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X439 a_22324_3994 a_21855_4398 VSS.t4 VSS.t3 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X440 VCTRL.t63 a_n17351_68.t37 EX.t29 VDD.t217 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X441 VSS.t257 a_24383_217 a_24335_261 VSS.t69 nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X442 a_n8659_n1230 a_n8537_93.t13 a_n8471_219.t4 VSS.t275 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X443 VSS.t293 a_23883_3430 a_23795_3522 VSS.t292 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X444 a_n17351_68.t1 FREERUN.t38 VSS.t202 VSS.t201 nfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
X445 EX.t15 FREERUN.t39 VCTRL.t1 VSS.t203 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X446 LF.t35 a_n17351_68.t38 VCTRL.t64 VSS.t228 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X447 OUT.t0 DOWN.t9 a_25265_6933 VSS.t105 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X448 VDD.t238 a_n8471_219.t11 a_10813_2840 VDD.t237 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X449 a_n9701_6193 a_16431_6193 VSS.t13 ppolyf_u r_width=0.8u r_length=0.13m
X450 VCTRL.t29 FREERUN.t40 LF.t1 VDD.t196 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X451 a_24443_4907 a_24355_4951 VSS.t51 VSS.t50 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X452 a_n558_2704.t0 a_11009_2840 a_14645_2840 VDD.t28 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X453 EX.t14 FREERUN.t41 VCTRL.t0 VSS.t212 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X454 a_25265_7733 a_24755_6933 OUT.t4 VDD.t257 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X455 EX.t22 a_n17351_68.t39 VCTRL.t44 VDD.t178 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X456 a_1712_13773 a_5840_14213 VSS.t0 ppolyf_u_1k r_width=1u r_length=20u
X457 a_n8537_n1530.t1 a_n8537_93.t14 a_21891_6933 VSS.t276 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X458 VCTRL.t45 a_n17351_68.t40 EX.t23 VDD.t179 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X459 VSS.t205 a_22203_n358.t20 a_22115_n302.t1 VSS.t199 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X460 VCTRL.t46 a_n17351_68.t41 EX.t24 VDD.t180 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
R0 VSS.n2700 VSS.n391 108707
R1 VSS.n1563 VSS.n1562 71567.2
R2 VSS.n2700 VSS.n2699 63487.1
R3 VSS.n1510 VSS.t277 44684.9
R4 VSS.n1678 VSS.n1677 41487.9
R5 VSS.n1679 VSS.n1566 41443.1
R6 VSS.n1510 VSS.n1006 40731.1
R7 VSS.n1565 VSS.n1564 38820.7
R8 VSS.n1511 VSS.n1510 38116.5
R9 VSS.n1562 VSS.n964 17415.5
R10 VSS.n1013 VSS.n964 13283.7
R11 VSS.n273 VSS.n131 12018.2
R12 VSS.n391 VSS.n390 11767.2
R13 VSS.n390 VSS.n295 11262.4
R14 VSS.n3239 VSS.n3238 10496.9
R15 VSS.n1679 VSS.n1678 8427.59
R16 VSS.n755 VSS.n23 8157.71
R17 VSS.n684 VSS.n45 8157.71
R18 VSS.n576 VSS.n67 8157.71
R19 VSS.n193 VSS.n89 8157.71
R20 VSS.n1510 VSS.n964 7822.41
R21 VSS.n2820 VSS.n194 7592.86
R22 VSS.n1866 VSS.n1837 7312.98
R23 VSS.n2413 VSS.n417 7297.55
R24 VSS.n3223 VSS.t296 6174.11
R25 VSS.n2595 VSS.n417 5958.33
R26 VSS.n275 VSS.n274 4966.24
R27 VSS.n2413 VSS.n2412 4966.24
R28 VSS.n3247 VSS.n3246 4888.01
R29 VSS.n1677 VSS.n1676 4674.55
R30 VSS.n1564 VSS.n1563 4034.48
R31 VSS.n277 VSS.n273 3373.39
R32 VSS.n3223 VSS.n131 2712.26
R33 VSS.n274 VSS.n98 2681.51
R34 VSS.t184 VSS.n118 2585.85
R35 VSS.n3246 VSS.n118 2574.44
R36 VSS.n329 VSS.n131 2530.6
R37 VSS.t13 VSS.n98 2437.5
R38 VSS.n3247 VSS.n111 2409.43
R39 VSS.n3229 VSS.n110 2232.27
R40 VSS.n3229 VSS.n118 2232.27
R41 VSS.n3255 VSS.n99 1975.11
R42 VSS.n3238 VSS.n3236 1861.31
R43 VSS.t233 VSS.t62 1662.1
R44 VSS.n1713 VSS.t210 1565.64
R45 VSS.n3236 VSS.n119 1540.41
R46 VSS.t199 VSS.t147 1513.7
R47 VSS.t13 VSS.n99 1503.17
R48 VSS.n274 VSS.n251 1460.46
R49 VSS.t71 VSS.t150 1439.5
R50 VSS.t206 VSS.n110 1421.85
R51 VSS.n1566 VSS.n1565 1412.07
R52 VSS.t81 VSS.t298 1406.11
R53 VSS.t60 VSS.t111 1394.98
R54 VSS.t113 VSS.t290 1365.3
R55 VSS.n410 VSS.t121 1362.36
R56 VSS.n1235 VSS.n1205 1310.22
R57 VSS.n1713 VSS.t138 1298.52
R58 VSS.t147 VSS.n1680 1261.42
R59 VSS.t79 VSS.t31 1250.29
R60 VSS.n1681 VSS.t71 1246.58
R61 VSS.n940 VSS.t210 1231.74
R62 VSS.t20 VSS.t242 1202.05
R63 VSS.t74 VSS.t35 1202.05
R64 VSS.n3188 VSS.t274 1191.86
R65 VSS.n3263 VSS.n3 1186.87
R66 VSS.n3263 VSS.n102 1171.01
R67 VSS.t5 VSS.t67 1157.53
R68 VSS.t56 VSS.n968 1113.01
R69 VSS.n962 VSS.t62 1113.01
R70 VSS.n967 VSS.t10 1109.3
R71 VSS.t288 VSS.t65 1101.88
R72 VSS.t9 VSS.t15 1101.88
R73 VSS.t231 VSS.t91 1044.49
R74 VSS.t179 VSS.t171 1044.49
R75 VSS.t150 VSS.t69 994.293
R76 VSS.n3253 VSS.n110 982.053
R77 VSS.t201 VSS.n111 982.053
R78 VSS.t250 VSS.t8 960.903
R79 VSS.n1633 VSS.t261 949.024
R80 VSS.n1944 VSS.t189 949.024
R81 VSS.n1978 VSS.t219 949.024
R82 VSS.n2221 VSS.t193 949.024
R83 VSS.n2255 VSS.t191 949.024
R84 VSS.n440 VSS.t259 949.024
R85 VSS.n330 VSS.n329 908.319
R86 VSS.n1564 VSS.n891 904.097
R87 VSS.n3223 VSS.t239 899.178
R88 VSS.t229 VSS.t175 889.111
R89 VSS.n1633 VSS.t216 873.673
R90 VSS.n1944 VSS.t40 873.673
R91 VSS.n1978 VSS.t249 873.673
R92 VSS.n2221 VSS.t58 873.673
R93 VSS.n2255 VSS.t120 873.673
R94 VSS.n440 VSS.t197 873.673
R95 VSS.n1837 VSS.n891 868.476
R96 VSS.t158 VSS.n963 845.89
R97 VSS.n970 VSS.n969 831.051
R98 VSS.t164 VSS.t73 831.051
R99 VSS.t73 VSS.t5 831.051
R100 VSS.t290 VSS.t199 831.051
R101 VSS.n3227 VSS.t268 782.889
R102 VSS.n3228 VSS.t245 769.885
R103 VSS.t7 VSS.t287 756.85
R104 VSS.t117 VSS.t263 756.85
R105 VSS.n1713 VSS.n934 749.429
R106 VSS.n1566 VSS.n912 728.482
R107 VSS.t263 VSS.t75 719.75
R108 VSS.n1563 VSS.n963 719.75
R109 VSS.n1565 VSS.n962 719.75
R110 VSS.n1680 VSS.n1679 719.75
R111 VSS.t11 VSS.t279 708.62
R112 VSS.t115 VSS.t11 686.359
R113 VSS.t118 VSS.t292 682.649
R114 VSS.t146 VSS.t115 682.649
R115 VSS.t279 VSS.t3 682.649
R116 VSS.t19 VSS.n943 682.649
R117 VSS.t235 VSS.t284 682.649
R118 VSS.t93 VSS.n1713 677.624
R119 VSS.n3224 VSS.n130 657.931
R120 VSS.t264 VSS.t48 649.259
R121 VSS.t171 VSS.n928 647.41
R122 VSS.t142 VSS.t46 638.129
R123 VSS.n945 VSS.t264 626.999
R124 VSS.t46 VSS.t103 623.288
R125 VSS.t69 VSS.t164 623.288
R126 VSS.t67 VSS.t74 623.288
R127 VSS.t35 VSS.t113 623.288
R128 VSS.n3206 VSS.n3204 617.557
R129 VSS.n2697 VSS.n394 583.484
R130 VSS.n2691 VSS.n394 583.484
R131 VSS.n2691 VSS.n2690 583.484
R132 VSS.n2690 VSS.n2689 583.484
R133 VSS.n2689 VSS.n2669 583.484
R134 VSS.n2683 VSS.n2669 583.484
R135 VSS.n2683 VSS.n2682 583.484
R136 VSS.n2682 VSS.n2681 583.484
R137 VSS.n2681 VSS.n2673 583.484
R138 VSS.n2675 VSS.n2673 583.484
R139 VSS.n2675 VSS.n124 583.484
R140 VSS.n3239 VSS.n124 583.484
R141 VSS.n2698 VSS.n2697 583.271
R142 VSS.t127 VSS.t33 567.638
R143 VSS.n251 VSS.n194 564.85
R144 VSS.t17 VSS.t288 560.217
R145 VSS.t165 VSS.n934 549.087
R146 VSS.t286 VSS.t255 549.087
R147 VSS.n968 VSS.t118 549.087
R148 VSS.n1675 VSS.n1571 534.539
R149 VSS.n1669 VSS.n1668 534.539
R150 VSS.n1668 VSS.n1667 534.539
R151 VSS.n1667 VSS.n1627 534.539
R152 VSS.n1661 VSS.n1627 534.539
R153 VSS.n1661 VSS.n1660 534.539
R154 VSS.n1660 VSS.n1659 534.539
R155 VSS.n1659 VSS.n1631 534.539
R156 VSS.n1652 VSS.n1631 534.539
R157 VSS.n1652 VSS.n1651 534.539
R158 VSS.n1651 VSS.n1650 534.539
R159 VSS.n1650 VSS.n1636 534.539
R160 VSS.n1644 VSS.n1636 534.539
R161 VSS.n1644 VSS.n1643 534.539
R162 VSS.n1643 VSS.n1642 534.539
R163 VSS.n1642 VSS.n811 534.539
R164 VSS.n1924 VSS.n811 534.539
R165 VSS.n1931 VSS.n1930 534.539
R166 VSS.n1932 VSS.n1931 534.539
R167 VSS.n1932 VSS.n802 534.539
R168 VSS.n1938 VSS.n802 534.539
R169 VSS.n1939 VSS.n1938 534.539
R170 VSS.n1940 VSS.n1939 534.539
R171 VSS.n1940 VSS.n798 534.539
R172 VSS.n1948 VSS.n798 534.539
R173 VSS.n1949 VSS.n1948 534.539
R174 VSS.n1950 VSS.n1949 534.539
R175 VSS.n1950 VSS.n794 534.539
R176 VSS.n1956 VSS.n794 534.539
R177 VSS.n1957 VSS.n1956 534.539
R178 VSS.n1958 VSS.n1957 534.539
R179 VSS.n1958 VSS.n790 534.539
R180 VSS.n1964 VSS.n790 534.539
R181 VSS.n1965 VSS.n1964 534.539
R182 VSS.n1966 VSS.n1965 534.539
R183 VSS.n2020 VSS.n2019 534.539
R184 VSS.n2019 VSS.n2018 534.539
R185 VSS.n2018 VSS.n1972 534.539
R186 VSS.n2012 VSS.n1972 534.539
R187 VSS.n2012 VSS.n2011 534.539
R188 VSS.n2011 VSS.n2010 534.539
R189 VSS.n2010 VSS.n1976 534.539
R190 VSS.n2004 VSS.n1976 534.539
R191 VSS.n2004 VSS.n2003 534.539
R192 VSS.n2003 VSS.n2002 534.539
R193 VSS.n2002 VSS.n1981 534.539
R194 VSS.n1996 VSS.n1981 534.539
R195 VSS.n1996 VSS.n1995 534.539
R196 VSS.n1995 VSS.n1994 534.539
R197 VSS.n1994 VSS.n1986 534.539
R198 VSS.n1988 VSS.n1986 534.539
R199 VSS.n1988 VSS.n632 534.539
R200 VSS.n2201 VSS.n632 534.539
R201 VSS.n2208 VSS.n2207 534.539
R202 VSS.n2209 VSS.n2208 534.539
R203 VSS.n2209 VSS.n623 534.539
R204 VSS.n2215 VSS.n623 534.539
R205 VSS.n2216 VSS.n2215 534.539
R206 VSS.n2217 VSS.n2216 534.539
R207 VSS.n2217 VSS.n619 534.539
R208 VSS.n2225 VSS.n619 534.539
R209 VSS.n2226 VSS.n2225 534.539
R210 VSS.n2227 VSS.n2226 534.539
R211 VSS.n2227 VSS.n615 534.539
R212 VSS.n2233 VSS.n615 534.539
R213 VSS.n2234 VSS.n2233 534.539
R214 VSS.n2235 VSS.n2234 534.539
R215 VSS.n2235 VSS.n611 534.539
R216 VSS.n2241 VSS.n611 534.539
R217 VSS.n2242 VSS.n2241 534.539
R218 VSS.n2243 VSS.n2242 534.539
R219 VSS.n2297 VSS.n2296 534.539
R220 VSS.n2296 VSS.n2295 534.539
R221 VSS.n2295 VSS.n2249 534.539
R222 VSS.n2289 VSS.n2249 534.539
R223 VSS.n2289 VSS.n2288 534.539
R224 VSS.n2288 VSS.n2287 534.539
R225 VSS.n2287 VSS.n2253 534.539
R226 VSS.n2281 VSS.n2253 534.539
R227 VSS.n2281 VSS.n2280 534.539
R228 VSS.n2280 VSS.n2279 534.539
R229 VSS.n2279 VSS.n2258 534.539
R230 VSS.n2273 VSS.n2258 534.539
R231 VSS.n2273 VSS.n2272 534.539
R232 VSS.n2272 VSS.n2271 534.539
R233 VSS.n2271 VSS.n2263 534.539
R234 VSS.n2265 VSS.n2263 534.539
R235 VSS.n2265 VSS.n453 534.539
R236 VSS.n2528 VSS.n453 534.539
R237 VSS.n2535 VSS.n447 534.539
R238 VSS.n2536 VSS.n2535 534.539
R239 VSS.n2537 VSS.n2536 534.539
R240 VSS.n2537 VSS.n443 534.539
R241 VSS.n2543 VSS.n443 534.539
R242 VSS.n2544 VSS.n2543 534.539
R243 VSS.n2545 VSS.n2544 534.539
R244 VSS.n2545 VSS.n438 534.539
R245 VSS.n2552 VSS.n438 534.539
R246 VSS.n2553 VSS.n2552 534.539
R247 VSS.n2554 VSS.n2553 534.539
R248 VSS.n2554 VSS.n434 534.539
R249 VSS.n2560 VSS.n434 534.539
R250 VSS.n2561 VSS.n2560 534.539
R251 VSS.n2563 VSS.n2561 534.539
R252 VSS.n2563 VSS.n2562 534.539
R253 VSS.n2562 VSS.n430 534.539
R254 VSS.n2586 VSS.n2585 534.539
R255 VSS.n2588 VSS.n2586 534.539
R256 VSS.n2588 VSS.n2587 534.539
R257 VSS.n3205 VSS.n129 533.557
R258 VSS.t25 VSS.t26 519.268
R259 VSS.t275 VSS.t25 519.268
R260 VSS.t268 VSS.t275 519.268
R261 VSS.t130 VSS.t160 510.158
R262 VSS.t136 VSS.t130 510.158
R263 VSS.t245 VSS.t136 510.158
R264 VSS.n1669 VSS.n1626 494.45
R265 VSS.t1 VSS.t265 486.017
R266 VSS.t144 VSS.n1555 484.224
R267 VSS.t95 VSS.t93 483.401
R268 VSS.t99 VSS.t95 483.401
R269 VSS.t87 VSS.t99 483.401
R270 VSS.t97 VSS.t87 483.401
R271 VSS.t101 VSS.t97 483.401
R272 VSS.t89 VSS.t101 483.401
R273 VSS.t91 VSS.t89 483.401
R274 VSS.t236 VSS.t229 483.401
R275 VSS.t175 VSS.t177 483.401
R276 VSS.t177 VSS.t173 483.401
R277 VSS.t173 VSS.t179 483.401
R278 VSS.t13 VSS.n100 444.149
R279 VSS.n3255 VSS.n3254 435.764
R280 VSS.t292 VSS.n967 430.365
R281 VSS.t77 VSS.t19 430.365
R282 VSS.n1677 VSS.n928 418.659
R283 VSS.n1236 VSS.n1081 416.675
R284 VSS.n1488 VSS.n1487 403.765
R285 VSS.n1487 VSS.n1486 403.765
R286 VSS.n1486 VSS.n1066 403.765
R287 VSS.n1480 VSS.n1066 403.765
R288 VSS.n1480 VSS.n1479 403.765
R289 VSS.n1479 VSS.n1478 403.765
R290 VSS.n1478 VSS.n1070 403.765
R291 VSS.t103 VSS.t77 400.685
R292 VSS.n1556 VSS.t132 394.5
R293 VSS.n1784 VSS.n916 388.524
R294 VSS.n1777 VSS.n890 388.524
R295 VSS.n1777 VSS.n1776 388.524
R296 VSS.n1776 VSS.n1775 388.524
R297 VSS.n1775 VSS.n1735 388.524
R298 VSS.n1769 VSS.n1735 388.524
R299 VSS.n1769 VSS.n1768 388.524
R300 VSS.n1768 VSS.n1767 388.524
R301 VSS.n1767 VSS.n1740 388.524
R302 VSS.n1761 VSS.n1740 388.524
R303 VSS.n1761 VSS.n1760 388.524
R304 VSS.n1760 VSS.n1759 388.524
R305 VSS.n1759 VSS.n1744 388.524
R306 VSS.n1753 VSS.n1744 388.524
R307 VSS.n1753 VSS.n1752 388.524
R308 VSS.n1752 VSS.n1751 388.524
R309 VSS.n1751 VSS.n828 388.524
R310 VSS.n885 VSS.n884 388.524
R311 VSS.n884 VSS.n883 388.524
R312 VSS.n883 VSS.n837 388.524
R313 VSS.n877 VSS.n837 388.524
R314 VSS.n877 VSS.n876 388.524
R315 VSS.n876 VSS.n875 388.524
R316 VSS.n875 VSS.n842 388.524
R317 VSS.n869 VSS.n842 388.524
R318 VSS.n869 VSS.n868 388.524
R319 VSS.n868 VSS.n867 388.524
R320 VSS.n867 VSS.n846 388.524
R321 VSS.n861 VSS.n846 388.524
R322 VSS.n861 VSS.n860 388.524
R323 VSS.n860 VSS.n859 388.524
R324 VSS.n859 VSS.n850 388.524
R325 VSS.n853 VSS.n850 388.524
R326 VSS.n853 VSS.n718 388.524
R327 VSS.n2062 VSS.n718 388.524
R328 VSS.n2067 VSS.n2066 388.524
R329 VSS.n2067 VSS.n711 388.524
R330 VSS.n2073 VSS.n711 388.524
R331 VSS.n2074 VSS.n2073 388.524
R332 VSS.n2075 VSS.n2074 388.524
R333 VSS.n2075 VSS.n707 388.524
R334 VSS.n2081 VSS.n707 388.524
R335 VSS.n2082 VSS.n2081 388.524
R336 VSS.n2083 VSS.n2082 388.524
R337 VSS.n2083 VSS.n703 388.524
R338 VSS.n2089 VSS.n703 388.524
R339 VSS.n2090 VSS.n2089 388.524
R340 VSS.n2091 VSS.n2090 388.524
R341 VSS.n2091 VSS.n699 388.524
R342 VSS.n2098 VSS.n699 388.524
R343 VSS.n2099 VSS.n2098 388.524
R344 VSS.n2100 VSS.n2099 388.524
R345 VSS.n2100 VSS.n649 388.524
R346 VSS.n2152 VSS.n2151 388.524
R347 VSS.n2151 VSS.n2150 388.524
R348 VSS.n2150 VSS.n2105 388.524
R349 VSS.n2144 VSS.n2105 388.524
R350 VSS.n2144 VSS.n2143 388.524
R351 VSS.n2143 VSS.n2142 388.524
R352 VSS.n2142 VSS.n2109 388.524
R353 VSS.n2136 VSS.n2109 388.524
R354 VSS.n2136 VSS.n2135 388.524
R355 VSS.n2135 VSS.n2134 388.524
R356 VSS.n2134 VSS.n2113 388.524
R357 VSS.n2128 VSS.n2113 388.524
R358 VSS.n2128 VSS.n2127 388.524
R359 VSS.n2127 VSS.n2126 388.524
R360 VSS.n2126 VSS.n2117 388.524
R361 VSS.n2120 VSS.n2117 388.524
R362 VSS.n2120 VSS.n539 388.524
R363 VSS.n2339 VSS.n539 388.524
R364 VSS.n2344 VSS.n2343 388.524
R365 VSS.n2344 VSS.n532 388.524
R366 VSS.n2350 VSS.n532 388.524
R367 VSS.n2351 VSS.n2350 388.524
R368 VSS.n2352 VSS.n2351 388.524
R369 VSS.n2352 VSS.n528 388.524
R370 VSS.n2358 VSS.n528 388.524
R371 VSS.n2359 VSS.n2358 388.524
R372 VSS.n2360 VSS.n2359 388.524
R373 VSS.n2360 VSS.n524 388.524
R374 VSS.n2366 VSS.n524 388.524
R375 VSS.n2367 VSS.n2366 388.524
R376 VSS.n2368 VSS.n2367 388.524
R377 VSS.n2368 VSS.n520 388.524
R378 VSS.n2375 VSS.n520 388.524
R379 VSS.n2376 VSS.n2375 388.524
R380 VSS.n2377 VSS.n2376 388.524
R381 VSS.n2377 VSS.n474 388.524
R382 VSS.n2481 VSS.n192 388.524
R383 VSS.n2481 VSS.n2480 388.524
R384 VSS.n2480 VSS.n2479 388.524
R385 VSS.n2479 VSS.n2383 388.524
R386 VSS.n2473 VSS.n2383 388.524
R387 VSS.n2473 VSS.n2472 388.524
R388 VSS.n2472 VSS.n2471 388.524
R389 VSS.n2471 VSS.n2388 388.524
R390 VSS.n2465 VSS.n2388 388.524
R391 VSS.n2465 VSS.n2464 388.524
R392 VSS.n2464 VSS.n2463 388.524
R393 VSS.n2463 VSS.n2392 388.524
R394 VSS.n2457 VSS.n2392 388.524
R395 VSS.n2457 VSS.n2456 388.524
R396 VSS.n2456 VSS.n2455 388.524
R397 VSS.n2455 VSS.n2396 388.524
R398 VSS.n2743 VSS.n2742 388.524
R399 VSS.n2742 VSS.n2741 388.524
R400 VSS.n2741 VSS.n265 388.524
R401 VSS.t296 VSS.t221 387.993
R402 VSS.t221 VSS.t167 387.993
R403 VSS.t167 VSS.t294 387.993
R404 VSS.t294 VSS.t183 387.993
R405 VSS.t183 VSS.t168 387.993
R406 VSS.t168 VSS.t181 387.993
R407 VSS.t181 VSS.t185 387.993
R408 VSS.t185 VSS.t186 387.993
R409 VSS.t186 VSS.t188 387.993
R410 VSS.t212 VSS.t295 387.993
R411 VSS.t170 VSS.t212 387.993
R412 VSS.t203 VSS.t170 387.993
R413 VSS.t169 VSS.t187 387.993
R414 VSS.t187 VSS.t182 387.993
R415 VSS.t182 VSS.t195 387.993
R416 VSS.t195 VSS.t153 387.993
R417 VSS.t153 VSS.t184 387.993
R418 VSS.n1081 VSS.n2 384.562
R419 VSS.n2571 VSS.n430 379.524
R420 VSS.n1590 VSS.n1586 372.921
R421 VSS.n1596 VSS.n1586 372.921
R422 VSS.n1597 VSS.n1596 372.921
R423 VSS.n1599 VSS.n1597 372.921
R424 VSS.n1599 VSS.n1598 372.921
R425 VSS.n1598 VSS.n1567 372.921
R426 VSS.n1581 VSS.n1568 372.921
R427 VSS.n1610 VSS.n1581 372.921
R428 VSS.n1611 VSS.n1610 372.921
R429 VSS.n1612 VSS.n1611 372.921
R430 VSS.n1612 VSS.n1576 372.921
R431 VSS.n1625 VSS.n1576 372.921
R432 VSS.n2587 VSS.n418 366.161
R433 VSS.n2412 VSS.n268 364.974
R434 VSS.n1224 VSS.t134 361.745
R435 VSS.t298 VSS.t142 356.164
R436 VSS.n384 VSS.n295 354.031
R437 VSS.n384 VSS.n383 354.031
R438 VSS.n383 VSS.n382 354.031
R439 VSS.n382 VSS.n132 354.031
R440 VSS.n3221 VSS.n132 354.031
R441 VSS.n1678 VSS.n1567 346.817
R442 VSS.n3222 VSS.n3221 341.639
R443 VSS.n1837 VSS.n889 336.074
R444 VSS.n3116 VSS.n99 332.938
R445 VSS.n1676 VSS.n1675 331.414
R446 VSS.n2585 VSS.n422 331.414
R447 VSS.n1714 VSS.t236 328.022
R448 VSS.n1626 VSS.n1625 324.442
R449 VSS.n2396 VSS.n194 316.647
R450 VSS.n2446 VSS.n2399 316.457
R451 VSS.n2440 VSS.n2439 316.457
R452 VSS.n2439 VSS.n2438 316.457
R453 VSS.n2438 VSS.n2414 316.457
R454 VSS.n2432 VSS.n2414 316.457
R455 VSS.n2430 VSS.n2429 316.457
R456 VSS.n2429 VSS.n2428 316.457
R457 VSS.n2428 VSS.n2418 316.457
R458 VSS.n2422 VSS.n2418 316.457
R459 VSS.n2572 VSS.n429 316.457
R460 VSS.n332 VSS.n330 310.856
R461 VSS.n1501 VSS.n1500 308.411
R462 VSS.n1502 VSS.n1501 308.411
R463 VSS.n1502 VSS.n1009 308.411
R464 VSS.n1508 VSS.n1009 308.411
R465 VSS.n1509 VSS.n1508 308.411
R466 VSS.n1511 VSS.n1509 308.411
R467 VSS.n1930 VSS.n806 307.361
R468 VSS.n2020 VSS.n1971 307.361
R469 VSS.n2207 VSS.n627 307.361
R470 VSS.n2297 VSS.n2248 307.361
R471 VSS.n2526 VSS.n447 307.361
R472 VSS.n1785 VSS.n912 306.935
R473 VSS.t54 VSS.t247 306.202
R474 VSS.n2597 VSS.n2596 302.748
R475 VSS.n2597 VSS.n413 302.748
R476 VSS.n2604 VSS.n413 302.748
R477 VSS.n2605 VSS.n2604 302.748
R478 VSS.n2606 VSS.n2605 302.748
R479 VSS.n2606 VSS.n408 302.748
R480 VSS.n2612 VSS.n408 302.748
R481 VSS.n2613 VSS.n2612 302.748
R482 VSS.n2614 VSS.n2613 302.748
R483 VSS.n2614 VSS.n404 302.748
R484 VSS.n2620 VSS.n404 302.748
R485 VSS.n2621 VSS.n2620 302.748
R486 VSS.n2652 VSS.n2621 302.748
R487 VSS.n2660 VSS.n398 302.748
R488 VSS.n2661 VSS.n2660 302.748
R489 VSS.n2662 VSS.n2661 302.748
R490 VSS.n2662 VSS.n392 302.748
R491 VSS.n2699 VSS.n392 296.693
R492 VSS.t65 VSS.t146 293.094
R493 VSS.n3236 VSS.t169 289.853
R494 VSS.n3224 VSS.n3223 288.923
R495 VSS.n1924 VSS.n1923 288.651
R496 VSS.n1966 VSS.n785 288.651
R497 VSS.n2201 VSS.n2200 288.651
R498 VSS.n2243 VSS.n606 288.651
R499 VSS.n2528 VSS.n2527 288.651
R500 VSS.n2570 VSS.n422 288.651
R501 VSS.n3234 VSS.n125 286.461
R502 VSS.n3200 VSS.n128 286.447
R503 VSS.n970 VSS.t165 281.964
R504 VSS.n274 VSS.n273 277.757
R505 VSS.n2707 VSS.n287 277.659
R506 VSS.n2701 VSS.n287 277.659
R507 VSS.n2629 VSS.n293 277.659
R508 VSS.n2629 VSS.n2622 277.659
R509 VSS.t227 VSS.t239 275.425
R510 VSS.t226 VSS.t227 275.425
R511 VSS.t213 VSS.t226 275.425
R512 VSS.t204 VSS.t213 275.425
R513 VSS.t215 VSS.t204 275.425
R514 VSS.t241 VSS.t215 275.425
R515 VSS.t228 VSS.t241 275.425
R516 VSS.t207 VSS.t228 275.425
R517 VSS.t196 VSS.t207 275.425
R518 VSS.t223 VSS.t300 275.425
R519 VSS.t300 VSS.t224 275.425
R520 VSS.t224 VSS.t225 275.425
R521 VSS.t225 VSS.t208 275.425
R522 VSS.t208 VSS.t222 275.425
R523 VSS.t222 VSS.t214 275.425
R524 VSS.t214 VSS.t240 275.425
R525 VSS.t240 VSS.t238 275.425
R526 VSS.t238 VSS.t206 275.425
R527 VSS.n2572 VSS.n2571 275.317
R528 VSS.n2430 VSS.n417 273.735
R529 VSS.n1488 VSS.n1013 272.236
R530 VSS.t3 VSS.t60 270.834
R531 VSS.n1889 VSS.n1888 270.495
R532 VSS.n1889 VSS.n824 270.495
R533 VSS.n1895 VSS.n824 270.495
R534 VSS.n1896 VSS.n1895 270.495
R535 VSS.n1897 VSS.n1896 270.495
R536 VSS.n1897 VSS.n820 270.495
R537 VSS.n1903 VSS.n820 270.495
R538 VSS.n1904 VSS.n1903 270.495
R539 VSS.n1905 VSS.n1904 270.495
R540 VSS.n1905 VSS.n816 270.495
R541 VSS.n1912 VSS.n816 270.495
R542 VSS.n1913 VSS.n1912 270.495
R543 VSS.n1914 VSS.n1913 270.495
R544 VSS.n2059 VSS.n723 270.495
R545 VSS.n2053 VSS.n723 270.495
R546 VSS.n2053 VSS.n2052 270.495
R547 VSS.n2052 VSS.n2051 270.495
R548 VSS.n2051 VSS.n774 270.495
R549 VSS.n2045 VSS.n774 270.495
R550 VSS.n2045 VSS.n2044 270.495
R551 VSS.n2044 VSS.n2043 270.495
R552 VSS.n2043 VSS.n778 270.495
R553 VSS.n2037 VSS.n778 270.495
R554 VSS.n2037 VSS.n2036 270.495
R555 VSS.n2036 VSS.n2035 270.495
R556 VSS.n2035 VSS.n782 270.495
R557 VSS.n2166 VSS.n2165 270.495
R558 VSS.n2166 VSS.n645 270.495
R559 VSS.n2172 VSS.n645 270.495
R560 VSS.n2173 VSS.n2172 270.495
R561 VSS.n2174 VSS.n2173 270.495
R562 VSS.n2174 VSS.n641 270.495
R563 VSS.n2180 VSS.n641 270.495
R564 VSS.n2181 VSS.n2180 270.495
R565 VSS.n2182 VSS.n2181 270.495
R566 VSS.n2182 VSS.n637 270.495
R567 VSS.n2189 VSS.n637 270.495
R568 VSS.n2190 VSS.n2189 270.495
R569 VSS.n2191 VSS.n2190 270.495
R570 VSS.n2336 VSS.n544 270.495
R571 VSS.n2330 VSS.n544 270.495
R572 VSS.n2330 VSS.n2329 270.495
R573 VSS.n2329 VSS.n2328 270.495
R574 VSS.n2328 VSS.n595 270.495
R575 VSS.n2322 VSS.n595 270.495
R576 VSS.n2322 VSS.n2321 270.495
R577 VSS.n2321 VSS.n2320 270.495
R578 VSS.n2320 VSS.n599 270.495
R579 VSS.n2314 VSS.n599 270.495
R580 VSS.n2314 VSS.n2313 270.495
R581 VSS.n2313 VSS.n2312 270.495
R582 VSS.n2312 VSS.n603 270.495
R583 VSS.n2496 VSS.n470 270.495
R584 VSS.n2497 VSS.n2496 270.495
R585 VSS.n2498 VSS.n2497 270.495
R586 VSS.n2498 VSS.n466 270.495
R587 VSS.n2504 VSS.n466 270.495
R588 VSS.n2505 VSS.n2504 270.495
R589 VSS.n2506 VSS.n2505 270.495
R590 VSS.n2506 VSS.n462 270.495
R591 VSS.n2512 VSS.n462 270.495
R592 VSS.n2513 VSS.n2512 270.495
R593 VSS.n2514 VSS.n2513 270.495
R594 VSS.n2514 VSS.n457 270.495
R595 VSS.n2525 VSS.n457 270.495
R596 VSS.t111 VSS.t158 267.123
R597 VSS.t15 VSS.t138 267.123
R598 VSS.n1785 VSS.n1784 264.197
R599 VSS.n2743 VSS.n259 264.197
R600 VSS.n2708 VSS.n2707 263.776
R601 VSS.n969 VSS.t7 255.994
R602 VSS.t50 VSS.t253 254.93
R603 VSS.n3234 VSS.n126 253.106
R604 VSS.n3200 VSS.n112 253.106
R605 VSS.n2449 VSS.n2448 252.541
R606 VSS.n3203 VSS.n3202 249.606
R607 VSS.n3202 VSS.n142 249.606
R608 VSS.n3254 VSS.n3253 245.012
R609 VSS.t85 VSS.t272 243.536
R610 VSS.n3222 VSS.n130 242.852
R611 VSS.n2412 VSS.n265 242.827
R612 VSS.t269 VSS.t141 242.113
R613 VSS.t303 VSS.t105 242.113
R614 VSS.t162 VSS.t303 242.113
R615 VSS.t253 VSS.t109 242.113
R616 VSS.t156 VSS.t244 242.113
R617 VSS.t247 VSS.t304 242.113
R618 VSS.t243 VSS.t85 242.113
R619 VSS.t157 VSS.t276 242.113
R620 VSS.t276 VSS.t83 242.113
R621 VSS.n2700 VSS.n293 240.175
R622 VSS.n885 VSS.n23 237
R623 VSS.n2066 VSS.n45 237
R624 VSS.n2152 VSS.n67 237
R625 VSS.n2343 VSS.n89 237
R626 VSS.n2820 VSS.n192 237
R627 VSS.n1914 VSS.n806 235.332
R628 VSS.n1971 VSS.n782 235.332
R629 VSS.n2191 VSS.n627 235.332
R630 VSS.n2248 VSS.n603 235.332
R631 VSS.n2526 VSS.n2525 235.332
R632 VSS.t140 VSS.t129 232.143
R633 VSS.n3248 VSS.n117 226.763
R634 VSS.n1236 VSS.n935 207.988
R635 VSS.n1500 VSS.n1013 207.945
R636 VSS.n2726 VSS.n2725 207.668
R637 VSS.n2725 VSS.n2724 207.668
R638 VSS.n2724 VSS.n278 207.668
R639 VSS.n2718 VSS.n278 207.668
R640 VSS.n2718 VSS.n2717 207.668
R641 VSS.n2717 VSS.n2716 207.668
R642 VSS.n2716 VSS.n282 207.668
R643 VSS.n2710 VSS.n282 207.668
R644 VSS.n2710 VSS.n2709 207.668
R645 VSS.n372 VSS.n300 207.668
R646 VSS.n373 VSS.n372 207.668
R647 VSS.n374 VSS.n373 207.668
R648 VSS.n374 VSS.n294 207.668
R649 VSS.t8 VSS.t1 196.632
R650 VSS.n1715 VSS.n932 195.534
R651 VSS.n3235 VSS.t188 193.996
R652 VSS.t295 VSS.n3235 193.996
R653 VSS.n391 VSS.n294 191.054
R654 VSS.t41 VSS.t140 189.417
R655 VSS.n2650 VSS.n398 187.704
R656 VSS.n1886 VSS.n828 186.492
R657 VSS.n2062 VSS.n2061 186.492
R658 VSS.n2163 VSS.n649 186.492
R659 VSS.n2339 VSS.n2338 186.492
R660 VSS.n2489 VSS.n474 186.492
R661 VSS.n2447 VSS.n259 186.492
R662 VSS.n1235 VSS.n1234 176.641
R663 VSS.n2422 VSS.n418 172.469
R664 VSS.t255 VSS.t117 170.662
R665 VSS.n2413 VSS.n2399 164.558
R666 VSS.n1713 VSS.t24 163.782
R667 VSS.t45 VSS.n1198 161.487
R668 VSS.n2595 VSS.n2594 158.944
R669 VSS.n1714 VSS.t231 155.379
R670 VSS.n2571 VSS.n2570 155.017
R671 VSS.t123 VSS.t243 152.388
R672 VSS.n2440 VSS.n2413 151.899
R673 VSS.n1556 VSS.t272 150.964
R674 VSS.t282 VSS.t157 149.541
R675 VSS.n943 VSS.t250 148.403
R676 VSS.t52 VSS.n1204 148.343
R677 VSS.n1201 VSS.t104 147.215
R678 VSS.t31 VSS.t235 144.692
R679 VSS.n429 VSS.n418 143.988
R680 VSS.n1210 VSS.t27 143.844
R681 VSS.n2596 VSS.n2595 143.805
R682 VSS.t59 VSS.n1084 141.207
R683 VSS.t109 VSS.t154 140.995
R684 VSS.n1225 VSS.t50 139.571
R685 VSS.t280 VSS.t156 138.147
R686 VSS.n3201 VSS.t196 137.713
R687 VSS.n3201 VSS.t223 137.713
R688 VSS.t265 VSS.t20 137.273
R689 VSS.n2448 VSS.n2447 135.983
R690 VSS.n3240 VSS.n123 135.464
R691 VSS.t287 VSS.t286 133.562
R692 VSS.n276 VSS.n275 131.869
R693 VSS.n945 VSS.t9 129.852
R694 VSS.n277 VSS.n276 129.792
R695 VSS.n332 VSS.n331 124.343
R696 VSS.n1209 VSS.t24 123.904
R697 VSS.n3248 VSS.n113 122.868
R698 VSS.n3230 VSS.n112 122.868
R699 VSS.n3230 VSS.n126 122.868
R700 VSS.t10 VSS.t17 122.433
R701 VSS.t141 VSS.n1209 118.209
R702 VSS.t75 VSS.t56 115.011
R703 VSS.t33 VSS.t79 115.011
R704 VSS.t134 VSS.t280 103.966
R705 VSS.n126 VSS.n117 103.895
R706 VSS.n3252 VSS.n112 103.895
R707 VSS.n3252 VSS.n113 103.895
R708 VSS.t154 VSS.t162 101.118
R709 VSS.n275 VSS.n268 99.9337
R710 VSS.n1100 VSS.n1094 99.1454
R711 VSS.n1190 VSS.n1100 99.1454
R712 VSS.n1190 VSS.n1189 99.1454
R713 VSS.n1189 VSS.n1188 99.1454
R714 VSS.n1178 VSS.n1177 99.1454
R715 VSS.n1171 VSS.n1121 99.1454
R716 VSS.n1171 VSS.n1170 99.1454
R717 VSS.n1494 VSS.n1018 99.1454
R718 VSS.t244 VSS.n1210 98.2696
R719 VSS.n3236 VSS.t203 98.1395
R720 VSS.n2594 VSS.n418 95.3661
R721 VSS.n313 VSS.n312 94.601
R722 VSS.n319 VSS.n312 94.601
R723 VSS.n320 VSS.n319 94.601
R724 VSS.n321 VSS.n320 94.601
R725 VSS.t132 VSS.t282 92.5728
R726 VSS.t304 VSS.t123 89.7244
R727 VSS.n2652 VSS.n2651 87.7974
R728 VSS.n1234 VSS.t270 85.2434
R729 VSS.n1715 VSS.n933 82.7755
R730 VSS.n1177 VSS.n1112 82.6213
R731 VSS.n3206 VSS.n3205 81.2783
R732 VSS.n2726 VSS.n277 77.8759
R733 VSS.n331 VSS.n286 77.8759
R734 VSS.n2651 VSS.n2650 75.6875
R735 VSS.n2449 VSS.n194 71.8774
R736 VSS.n1170 VSS.n1017 69.8526
R737 VSS.n1198 VSS.n1094 65.346
R738 VSS.n3223 VSS.n3222 64.4305
R739 VSS.n3429 VSS.n2 63.438
R740 VSS.n331 VSS.n300 63.3392
R741 VSS.n1552 VSS.n992 62.7954
R742 VSS.n993 VSS.n964 60.9861
R743 VSS.n2651 VSS.n2622 59.6972
R744 VSS.t242 VSS.t127 55.6512
R745 VSS.n1517 VSS.n1516 54.8952
R746 VSS.n1156 VSS.n1155 53.1452
R747 VSS.n1816 VSS.n892 53.0314
R748 VSS.n1836 VSS.n893 53.0314
R749 VSS.n1830 VSS.n893 53.0314
R750 VSS.n1830 VSS.n1829 53.0314
R751 VSS.n1829 VSS.n1828 53.0314
R752 VSS.n1828 VSS.n1822 53.0314
R753 VSS.n1822 VSS.n4 53.0314
R754 VSS.n12 VSS.n5 53.0314
R755 VSS.n3419 VSS.n12 53.0314
R756 VSS.n3419 VSS.n3418 53.0314
R757 VSS.n3418 VSS.n3417 53.0314
R758 VSS.n3417 VSS.n13 53.0314
R759 VSS.n3411 VSS.n13 53.0314
R760 VSS.n3411 VSS.n3410 53.0314
R761 VSS.n3410 VSS.n3409 53.0314
R762 VSS.n3409 VSS.n17 53.0314
R763 VSS.n3402 VSS.n3401 53.0314
R764 VSS.n3401 VSS.n3400 53.0314
R765 VSS.n3400 VSS.n24 53.0314
R766 VSS.n3394 VSS.n24 53.0314
R767 VSS.n3394 VSS.n3393 53.0314
R768 VSS.n3393 VSS.n3392 53.0314
R769 VSS.n3392 VSS.n28 53.0314
R770 VSS.n3386 VSS.n28 53.0314
R771 VSS.n3386 VSS.n3385 53.0314
R772 VSS.n3385 VSS.n3384 53.0314
R773 VSS.n3384 VSS.n32 53.0314
R774 VSS.n3378 VSS.n32 53.0314
R775 VSS.n3378 VSS.n3377 53.0314
R776 VSS.n3377 VSS.n3376 53.0314
R777 VSS.n3376 VSS.n36 53.0314
R778 VSS.n3370 VSS.n36 53.0314
R779 VSS.n3370 VSS.n3369 53.0314
R780 VSS.n3369 VSS.n3368 53.0314
R781 VSS.n3362 VSS.n3361 53.0314
R782 VSS.n3361 VSS.n3360 53.0314
R783 VSS.n3360 VSS.n46 53.0314
R784 VSS.n3354 VSS.n46 53.0314
R785 VSS.n3354 VSS.n3353 53.0314
R786 VSS.n3353 VSS.n3352 53.0314
R787 VSS.n3352 VSS.n50 53.0314
R788 VSS.n3346 VSS.n50 53.0314
R789 VSS.n3346 VSS.n3345 53.0314
R790 VSS.n3345 VSS.n3344 53.0314
R791 VSS.n3344 VSS.n54 53.0314
R792 VSS.n3338 VSS.n54 53.0314
R793 VSS.n3338 VSS.n3337 53.0314
R794 VSS.n3337 VSS.n3336 53.0314
R795 VSS.n3336 VSS.n58 53.0314
R796 VSS.n3330 VSS.n58 53.0314
R797 VSS.n3330 VSS.n3329 53.0314
R798 VSS.n3329 VSS.n3328 53.0314
R799 VSS.n3322 VSS.n3321 53.0314
R800 VSS.n3321 VSS.n3320 53.0314
R801 VSS.n3320 VSS.n68 53.0314
R802 VSS.n3314 VSS.n68 53.0314
R803 VSS.n3314 VSS.n3313 53.0314
R804 VSS.n3313 VSS.n3312 53.0314
R805 VSS.n3312 VSS.n72 53.0314
R806 VSS.n3306 VSS.n72 53.0314
R807 VSS.n3306 VSS.n3305 53.0314
R808 VSS.n3305 VSS.n3304 53.0314
R809 VSS.n3304 VSS.n76 53.0314
R810 VSS.n3298 VSS.n76 53.0314
R811 VSS.n3298 VSS.n3297 53.0314
R812 VSS.n3297 VSS.n3296 53.0314
R813 VSS.n3296 VSS.n80 53.0314
R814 VSS.n3290 VSS.n80 53.0314
R815 VSS.n3290 VSS.n3289 53.0314
R816 VSS.n3289 VSS.n3288 53.0314
R817 VSS.n3282 VSS.n3281 53.0314
R818 VSS.n3281 VSS.n3280 53.0314
R819 VSS.n3280 VSS.n90 53.0314
R820 VSS.n3274 VSS.n90 53.0314
R821 VSS.n3274 VSS.n3273 53.0314
R822 VSS.n3273 VSS.n3272 53.0314
R823 VSS.n3266 VSS.n97 53.0314
R824 VSS.n208 VSS.n101 53.0314
R825 VSS.n209 VSS.n208 53.0314
R826 VSS.n210 VSS.n209 53.0314
R827 VSS.n210 VSS.n200 53.0314
R828 VSS.n217 VSS.n200 53.0314
R829 VSS.n218 VSS.n217 53.0314
R830 VSS.n219 VSS.n218 53.0314
R831 VSS.n219 VSS.n188 53.0314
R832 VSS.n2819 VSS.n195 53.0314
R833 VSS.n2813 VSS.n195 53.0314
R834 VSS.n2813 VSS.n2812 53.0314
R835 VSS.n2812 VSS.n2811 53.0314
R836 VSS.n2811 VSS.n226 53.0314
R837 VSS.n2805 VSS.n226 53.0314
R838 VSS.n2805 VSS.n2804 53.0314
R839 VSS.n2804 VSS.n2803 53.0314
R840 VSS.n2803 VSS.n230 53.0314
R841 VSS.n2797 VSS.n230 53.0314
R842 VSS.n2796 VSS.n2795 53.0314
R843 VSS.n2795 VSS.n234 53.0314
R844 VSS.n2789 VSS.n234 53.0314
R845 VSS.n2789 VSS.n2788 53.0314
R846 VSS.n2788 VSS.n2787 53.0314
R847 VSS.n2781 VSS.n241 53.0314
R848 VSS.n2779 VSS.n2773 53.0314
R849 VSS.n2773 VSS.n164 53.0314
R850 VSS.n3117 VSS.n164 53.0314
R851 VSS.n1196 VSS.n1195 52.7768
R852 VSS.n3264 VSS.n101 52.7663
R853 VSS.t105 VSS.t41 52.6955
R854 VSS.t270 VSS.t125 52.3156
R855 VSS.t125 VSS.t29 52.3156
R856 VSS.t29 VSS.t267 52.3156
R857 VSS.t23 VSS.t21 52.3156
R858 VSS.t22 VSS.t23 52.3156
R859 VSS.n1070 VSS.n964 52.0005
R860 VSS.n2708 VSS.n286 51.9174
R861 VSS.n313 VSS.n100 51.0848
R862 VSS.n1223 VSS.n935 50.2036
R863 VSS.n1837 VSS.n892 49.8496
R864 VSS.n1555 VSS.t277 49.8471
R865 VSS.n2709 VSS.n2708 47.7641
R866 VSS.n1837 VSS.n890 46.6233
R867 VSS.n2787 VSS.n194 46.4026
R868 VSS.n2432 VSS.n417 42.722
R869 VSS.n3266 VSS.t13 42.4252
R870 VSS.n1180 VSS.n1179 40.5598
R871 VSS.n1626 VSS.n1571 40.091
R872 VSS.n3272 VSS.t0 40.0388
R873 VSS.n1732 VSS.n919 39.3485
R874 VSS.n1573 VSS.n919 39.3305
R875 VSS.n3190 VSS.n111 38.8471
R876 VSS.t21 VSS.n1712 38.4675
R877 VSS.n3428 VSS.n4 38.4479
R878 VSS.n3253 VSS.t201 37.9805
R879 VSS.n2701 VSS.n2700 37.4845
R880 VSS.n1033 VSS.n1016 37.0268
R881 VSS.n2797 VSS.t14 36.857
R882 VSS.n3205 VSS.n128 36.8426
R883 VSS.n1061 VSS.n1019 36.6584
R884 VSS.n1550 VSS.n993 36.0615
R885 VSS.n3192 VSS.n3191 35.6452
R886 VSS.n3192 VSS.n112 35.6452
R887 VSS.n3191 VSS.n3190 35.6452
R888 VSS.n3190 VSS.n113 35.6452
R889 VSS.t38 VSS.n1104 33.4243
R890 VSS.n1183 VSS.t36 33.4243
R891 VSS.t48 VSS.t81 33.3909
R892 VSS.n1816 VSS.n1815 32.8797
R893 VSS.n2780 VSS.n2779 32.8797
R894 VSS.n1225 VSS.n1224 32.7569
R895 VSS.n1018 VSS.n1013 32.2977
R896 VSS.n1188 VSS.n1104 31.9222
R897 VSS.n1549 VSS.n1002 30.5794
R898 VSS.n3237 VSS.n123 30.2813
R899 VSS.n904 VSS.n896 29.7905
R900 VSS.n1732 VSS.n904 29.7725
R901 VSS.n1681 VSS.n940 29.6809
R902 VSS.n1494 VSS.n1017 29.2933
R903 VSS.n3402 VSS.n23 29.1675
R904 VSS.n3362 VSS.n45 29.1675
R905 VSS.n3322 VSS.n67 29.1675
R906 VSS.n3282 VSS.n89 29.1675
R907 VSS.n2820 VSS.n2819 29.1675
R908 VSS.n1847 VSS.n17 28.6372
R909 VSS.n3368 VSS.n40 28.6372
R910 VSS.n3328 VSS.n62 28.6372
R911 VSS.n3288 VSS.n84 28.6372
R912 VSS.n2781 VSS.n2780 28.6372
R913 VSS.n1545 VSS.n1544 28.3689
R914 VSS.n1541 VSS.n1540 28.3689
R915 VSS.n1537 VSS.n1536 28.3689
R916 VSS.n1533 VSS.n1532 28.3689
R917 VSS.n1529 VSS.n1528 28.3689
R918 VSS.n1525 VSS.n1524 28.3689
R919 VSS.n1521 VSS.n1520 28.3689
R920 VSS.n1061 VSS.n1060 28.0005
R921 VSS.n1058 VSS.n1022 28.0005
R922 VSS.n1054 VSS.n1053 28.0005
R923 VSS.n1051 VSS.n1025 28.0005
R924 VSS.n1047 VSS.n1046 28.0005
R925 VSS.n1044 VSS.n1028 28.0005
R926 VSS.n1040 VSS.n1039 28.0005
R927 VSS.n1037 VSS.n1031 28.0005
R928 VSS.n1096 VSS.n1095 28.0005
R929 VSS.n1126 VSS.n1095 28.0005
R930 VSS.n1130 VSS.n1129 28.0005
R931 VSS.n1134 VSS.n1133 28.0005
R932 VSS.n1138 VSS.n1137 28.0005
R933 VSS.n1142 VSS.n1141 28.0005
R934 VSS.n1146 VSS.n1145 28.0005
R935 VSS.n1150 VSS.n1149 28.0005
R936 VSS.n3245 VSS.n119 27.5094
R937 VSS.n1184 VSS.n1106 26.6645
R938 VSS.n1678 VSS.n1568 26.1049
R939 VSS.n1157 VSS.n1156 24.3163
R940 VSS.n1157 VSS.n1101 24.3163
R941 VSS.n1102 VSS.n1101 24.3163
R942 VSS.n1103 VSS.n1102 24.3163
R943 VSS.n1107 VSS.n1103 24.3163
R944 VSS.n1110 VSS.n1107 24.3163
R945 VSS.n1111 VSS.n1110 24.3163
R946 VSS.n1165 VSS.n1111 24.3163
R947 VSS.n1165 VSS.n1122 24.3163
R948 VSS.n1169 VSS.n1122 24.3163
R949 VSS.n1495 VSS.n1014 24.3163
R950 VSS.n1499 VSS.n1014 24.3163
R951 VSS.n1499 VSS.n1012 24.3163
R952 VSS.n1503 VSS.n1012 24.3163
R953 VSS.n1503 VSS.n1010 24.3163
R954 VSS.n1507 VSS.n1010 24.3163
R955 VSS.n1507 VSS.n1008 24.3163
R956 VSS.n1512 VSS.n1008 24.3163
R957 VSS.n1512 VSS.n1006 24.3163
R958 VSS.n1516 VSS.n1006 24.3163
R959 VSS.n1195 VSS.n1097 24.3163
R960 VSS.n1191 VSS.n1097 24.3163
R961 VSS.n1191 VSS.n1099 24.3163
R962 VSS.n1187 VSS.n1099 24.3163
R963 VSS.n1185 VSS.n1105 24.3163
R964 VSS.n1176 VSS.n1105 24.3163
R965 VSS.n1176 VSS.n1113 24.3163
R966 VSS.n1172 VSS.n1113 24.3163
R967 VSS.n1172 VSS.n1120 24.3163
R968 VSS.n1493 VSS.n1020 24.3163
R969 VSS.n1489 VSS.n1020 24.3163
R970 VSS.n1489 VSS.n1065 24.3163
R971 VSS.n1485 VSS.n1065 24.3163
R972 VSS.n1485 VSS.n1067 24.3163
R973 VSS.n1481 VSS.n1067 24.3163
R974 VSS.n1481 VSS.n1069 24.3163
R975 VSS.n1477 VSS.n1069 24.3163
R976 VSS.n1477 VSS.n1071 24.3163
R977 VSS.n1071 VSS.n1002 24.3163
R978 VSS.n1549 VSS.n1003 24.2242
R979 VSS.n1560 VSS.t278 24.116
R980 VSS.n1923 VSS.n806 24.0548
R981 VSS.n1971 VSS.n785 24.0548
R982 VSS.n2200 VSS.n627 24.0548
R983 VSS.n2248 VSS.n606 24.0548
R984 VSS.n2527 VSS.n2526 24.0548
R985 VSS.n1226 VSS.n1225 23.9005
R986 VSS.n1557 VSS.n1556 23.9005
R987 VSS.n1866 VSS.n23 23.7479
R988 VSS.n755 VSS.n45 23.7479
R989 VSS.n684 VSS.n67 23.7479
R990 VSS.n576 VSS.n89 23.7479
R991 VSS.n2820 VSS.n193 23.7479
R992 VSS.n1559 VSS.t84 22.3205
R993 VSS.n1558 VSS.t133 22.3205
R994 VSS.n965 VSS.t86 22.3205
R995 VSS.n1208 VSS.t135 22.3205
R996 VSS.n1227 VSS.t254 22.3205
R997 VSS.n1232 VSS.t271 22.3205
R998 VSS.n1551 VSS.n898 21.2129
R999 VSS.n1815 VSS.n898 20.6826
R1000 VSS.n1207 VSS.n1206 19.8005
R1001 VSS.n1229 VSS.n1228 19.8005
R1002 VSS.n1231 VSS.n1230 19.8005
R1003 VSS.n321 VSS.n131 18.9206
R1004 VSS.n247 VSS.n243 18.4216
R1005 VSS.n2771 VSS.n244 18.4216
R1006 VSS.n2767 VSS.n244 18.4216
R1007 VSS.n2765 VSS.n2764 18.4216
R1008 VSS.n2762 VSS.n253 18.4216
R1009 VSS.n2758 VSS.n2757 18.4216
R1010 VSS.n2755 VSS.n256 18.4216
R1011 VSS.n2751 VSS.n2750 18.4216
R1012 VSS.n488 VSS.n487 18.4216
R1013 VSS.n492 VSS.n491 18.4216
R1014 VSS.n494 VSS.n492 18.4216
R1015 VSS.n498 VSS.n482 18.4216
R1016 VSS.n502 VSS.n500 18.4216
R1017 VSS.n506 VSS.n480 18.4216
R1018 VSS.n509 VSS.n508 18.4216
R1019 VSS.n511 VSS.n477 18.4216
R1020 VSS.n559 VSS.n557 18.4216
R1021 VSS.n575 VSS.n552 18.4216
R1022 VSS.n575 VSS.n553 18.4216
R1023 VSS.n571 VSS.n570 18.4216
R1024 VSS.n567 VSS.n566 18.4216
R1025 VSS.n563 VSS.n548 18.4216
R1026 VSS.n579 VSS.n578 18.4216
R1027 VSS.n583 VSS.n582 18.4216
R1028 VSS.n1880 VSS.n832 18.4216
R1029 VSS.n1884 VSS.n827 18.4216
R1030 VSS.n1890 VSS.n827 18.4216
R1031 VSS.n1890 VSS.n825 18.4216
R1032 VSS.n1894 VSS.n825 18.4216
R1033 VSS.n1894 VSS.n823 18.4216
R1034 VSS.n1898 VSS.n823 18.4216
R1035 VSS.n1898 VSS.n821 18.4216
R1036 VSS.n1902 VSS.n821 18.4216
R1037 VSS.n1902 VSS.n819 18.4216
R1038 VSS.n1906 VSS.n819 18.4216
R1039 VSS.n1906 VSS.n817 18.4216
R1040 VSS.n1911 VSS.n817 18.4216
R1041 VSS.n1911 VSS.n815 18.4216
R1042 VSS.n1915 VSS.n815 18.4216
R1043 VSS.n1916 VSS.n1915 18.4216
R1044 VSS.n1920 VSS.n813 18.4216
R1045 VSS.n769 VSS.n768 18.4216
R1046 VSS.n2058 VSS.n724 18.4216
R1047 VSS.n2058 VSS.n725 18.4216
R1048 VSS.n2054 VSS.n725 18.4216
R1049 VSS.n2054 VSS.n773 18.4216
R1050 VSS.n2050 VSS.n773 18.4216
R1051 VSS.n2050 VSS.n775 18.4216
R1052 VSS.n2046 VSS.n775 18.4216
R1053 VSS.n2046 VSS.n777 18.4216
R1054 VSS.n2042 VSS.n777 18.4216
R1055 VSS.n2042 VSS.n779 18.4216
R1056 VSS.n2038 VSS.n779 18.4216
R1057 VSS.n2038 VSS.n781 18.4216
R1058 VSS.n2034 VSS.n781 18.4216
R1059 VSS.n2034 VSS.n783 18.4216
R1060 VSS.n2030 VSS.n783 18.4216
R1061 VSS.n2028 VSS.n2027 18.4216
R1062 VSS.n2161 VSS.n654 18.4216
R1063 VSS.n2157 VSS.n648 18.4216
R1064 VSS.n2167 VSS.n648 18.4216
R1065 VSS.n2167 VSS.n646 18.4216
R1066 VSS.n2171 VSS.n646 18.4216
R1067 VSS.n2171 VSS.n644 18.4216
R1068 VSS.n2175 VSS.n644 18.4216
R1069 VSS.n2175 VSS.n642 18.4216
R1070 VSS.n2179 VSS.n642 18.4216
R1071 VSS.n2179 VSS.n640 18.4216
R1072 VSS.n2183 VSS.n640 18.4216
R1073 VSS.n2183 VSS.n638 18.4216
R1074 VSS.n2188 VSS.n638 18.4216
R1075 VSS.n2188 VSS.n636 18.4216
R1076 VSS.n2192 VSS.n636 18.4216
R1077 VSS.n2193 VSS.n2192 18.4216
R1078 VSS.n2197 VSS.n634 18.4216
R1079 VSS.n590 VSS.n589 18.4216
R1080 VSS.n2335 VSS.n545 18.4216
R1081 VSS.n2335 VSS.n546 18.4216
R1082 VSS.n2331 VSS.n546 18.4216
R1083 VSS.n2331 VSS.n594 18.4216
R1084 VSS.n2327 VSS.n594 18.4216
R1085 VSS.n2327 VSS.n596 18.4216
R1086 VSS.n2323 VSS.n596 18.4216
R1087 VSS.n2323 VSS.n598 18.4216
R1088 VSS.n2319 VSS.n598 18.4216
R1089 VSS.n2319 VSS.n600 18.4216
R1090 VSS.n2315 VSS.n600 18.4216
R1091 VSS.n2315 VSS.n602 18.4216
R1092 VSS.n2311 VSS.n602 18.4216
R1093 VSS.n2311 VSS.n604 18.4216
R1094 VSS.n2307 VSS.n604 18.4216
R1095 VSS.n2305 VSS.n2304 18.4216
R1096 VSS.n514 VSS.n473 18.4216
R1097 VSS.n2491 VSS.n471 18.4216
R1098 VSS.n2495 VSS.n471 18.4216
R1099 VSS.n2495 VSS.n469 18.4216
R1100 VSS.n2499 VSS.n469 18.4216
R1101 VSS.n2499 VSS.n467 18.4216
R1102 VSS.n2503 VSS.n467 18.4216
R1103 VSS.n2503 VSS.n465 18.4216
R1104 VSS.n2507 VSS.n465 18.4216
R1105 VSS.n2507 VSS.n463 18.4216
R1106 VSS.n2511 VSS.n463 18.4216
R1107 VSS.n2511 VSS.n461 18.4216
R1108 VSS.n2515 VSS.n461 18.4216
R1109 VSS.n2515 VSS.n458 18.4216
R1110 VSS.n2524 VSS.n458 18.4216
R1111 VSS.n2524 VSS.n459 18.4216
R1112 VSS.n2520 VSS.n2519 18.4216
R1113 VSS.n667 VSS.n665 18.4216
R1114 VSS.n683 VSS.n660 18.4216
R1115 VSS.n683 VSS.n661 18.4216
R1116 VSS.n679 VSS.n678 18.4216
R1117 VSS.n675 VSS.n674 18.4216
R1118 VSS.n671 VSS.n656 18.4216
R1119 VSS.n687 VSS.n686 18.4216
R1120 VSS.n691 VSS.n690 18.4216
R1121 VSS.n2407 VSS.n2405 18.4216
R1122 VSS.n2445 VSS.n2400 18.4216
R1123 VSS.n2445 VSS.n2401 18.4216
R1124 VSS.n2441 VSS.n2401 18.4216
R1125 VSS.n2441 VSS.n2411 18.4216
R1126 VSS.n2437 VSS.n2411 18.4216
R1127 VSS.n2437 VSS.n2415 18.4216
R1128 VSS.n2433 VSS.n2415 18.4216
R1129 VSS.n2433 VSS.n2431 18.4216
R1130 VSS.n2431 VSS.n2417 18.4216
R1131 VSS.n2427 VSS.n2417 18.4216
R1132 VSS.n2427 VSS.n2419 18.4216
R1133 VSS.n2423 VSS.n2419 18.4216
R1134 VSS.n2423 VSS.n428 18.4216
R1135 VSS.n2573 VSS.n428 18.4216
R1136 VSS.n2574 VSS.n2573 18.4216
R1137 VSS.n2578 VSS.n2577 18.4216
R1138 VSS.n1674 VSS.n1572 18.4216
R1139 VSS.n1670 VSS.n1572 18.4216
R1140 VSS.n1670 VSS.n1575 18.4216
R1141 VSS.n1666 VSS.n1575 18.4216
R1142 VSS.n1666 VSS.n1628 18.4216
R1143 VSS.n1662 VSS.n1628 18.4216
R1144 VSS.n1662 VSS.n1630 18.4216
R1145 VSS.n1658 VSS.n1630 18.4216
R1146 VSS.n1658 VSS.n1632 18.4216
R1147 VSS.n1653 VSS.n1632 18.4216
R1148 VSS.n1653 VSS.n1635 18.4216
R1149 VSS.n1649 VSS.n1635 18.4216
R1150 VSS.n1649 VSS.n1637 18.4216
R1151 VSS.n1645 VSS.n1637 18.4216
R1152 VSS.n1645 VSS.n1639 18.4216
R1153 VSS.n1641 VSS.n1639 18.4216
R1154 VSS.n1641 VSS.n810 18.4216
R1155 VSS.n1925 VSS.n810 18.4216
R1156 VSS.n1929 VSS.n805 18.4216
R1157 VSS.n1933 VSS.n805 18.4216
R1158 VSS.n1933 VSS.n803 18.4216
R1159 VSS.n1937 VSS.n803 18.4216
R1160 VSS.n1937 VSS.n801 18.4216
R1161 VSS.n1941 VSS.n801 18.4216
R1162 VSS.n1941 VSS.n799 18.4216
R1163 VSS.n1947 VSS.n799 18.4216
R1164 VSS.n1947 VSS.n797 18.4216
R1165 VSS.n1951 VSS.n797 18.4216
R1166 VSS.n1951 VSS.n795 18.4216
R1167 VSS.n1955 VSS.n795 18.4216
R1168 VSS.n1955 VSS.n793 18.4216
R1169 VSS.n1959 VSS.n793 18.4216
R1170 VSS.n1959 VSS.n791 18.4216
R1171 VSS.n1963 VSS.n791 18.4216
R1172 VSS.n1963 VSS.n789 18.4216
R1173 VSS.n1967 VSS.n789 18.4216
R1174 VSS.n2021 VSS.n1970 18.4216
R1175 VSS.n2017 VSS.n1970 18.4216
R1176 VSS.n2017 VSS.n1973 18.4216
R1177 VSS.n2013 VSS.n1973 18.4216
R1178 VSS.n2013 VSS.n1975 18.4216
R1179 VSS.n2009 VSS.n1975 18.4216
R1180 VSS.n2009 VSS.n1977 18.4216
R1181 VSS.n2005 VSS.n1977 18.4216
R1182 VSS.n2005 VSS.n1980 18.4216
R1183 VSS.n2001 VSS.n1980 18.4216
R1184 VSS.n2001 VSS.n1982 18.4216
R1185 VSS.n1997 VSS.n1982 18.4216
R1186 VSS.n1997 VSS.n1985 18.4216
R1187 VSS.n1993 VSS.n1985 18.4216
R1188 VSS.n1993 VSS.n1987 18.4216
R1189 VSS.n1989 VSS.n1987 18.4216
R1190 VSS.n1989 VSS.n631 18.4216
R1191 VSS.n2202 VSS.n631 18.4216
R1192 VSS.n2206 VSS.n626 18.4216
R1193 VSS.n2210 VSS.n626 18.4216
R1194 VSS.n2210 VSS.n624 18.4216
R1195 VSS.n2214 VSS.n624 18.4216
R1196 VSS.n2214 VSS.n622 18.4216
R1197 VSS.n2218 VSS.n622 18.4216
R1198 VSS.n2218 VSS.n620 18.4216
R1199 VSS.n2224 VSS.n620 18.4216
R1200 VSS.n2224 VSS.n618 18.4216
R1201 VSS.n2228 VSS.n618 18.4216
R1202 VSS.n2228 VSS.n616 18.4216
R1203 VSS.n2232 VSS.n616 18.4216
R1204 VSS.n2232 VSS.n614 18.4216
R1205 VSS.n2236 VSS.n614 18.4216
R1206 VSS.n2236 VSS.n612 18.4216
R1207 VSS.n2240 VSS.n612 18.4216
R1208 VSS.n2240 VSS.n610 18.4216
R1209 VSS.n2244 VSS.n610 18.4216
R1210 VSS.n2298 VSS.n2247 18.4216
R1211 VSS.n2294 VSS.n2247 18.4216
R1212 VSS.n2294 VSS.n2250 18.4216
R1213 VSS.n2290 VSS.n2250 18.4216
R1214 VSS.n2290 VSS.n2252 18.4216
R1215 VSS.n2286 VSS.n2252 18.4216
R1216 VSS.n2286 VSS.n2254 18.4216
R1217 VSS.n2282 VSS.n2254 18.4216
R1218 VSS.n2282 VSS.n2257 18.4216
R1219 VSS.n2278 VSS.n2257 18.4216
R1220 VSS.n2278 VSS.n2259 18.4216
R1221 VSS.n2274 VSS.n2259 18.4216
R1222 VSS.n2274 VSS.n2262 18.4216
R1223 VSS.n2270 VSS.n2262 18.4216
R1224 VSS.n2270 VSS.n2264 18.4216
R1225 VSS.n2266 VSS.n2264 18.4216
R1226 VSS.n2266 VSS.n451 18.4216
R1227 VSS.n2529 VSS.n451 18.4216
R1228 VSS.n2534 VSS.n448 18.4216
R1229 VSS.n2534 VSS.n446 18.4216
R1230 VSS.n2538 VSS.n446 18.4216
R1231 VSS.n2538 VSS.n444 18.4216
R1232 VSS.n2542 VSS.n444 18.4216
R1233 VSS.n2542 VSS.n442 18.4216
R1234 VSS.n2546 VSS.n442 18.4216
R1235 VSS.n2546 VSS.n439 18.4216
R1236 VSS.n2551 VSS.n439 18.4216
R1237 VSS.n2551 VSS.n437 18.4216
R1238 VSS.n2555 VSS.n437 18.4216
R1239 VSS.n2555 VSS.n435 18.4216
R1240 VSS.n2559 VSS.n435 18.4216
R1241 VSS.n2559 VSS.n433 18.4216
R1242 VSS.n2564 VSS.n433 18.4216
R1243 VSS.n2564 VSS.n431 18.4216
R1244 VSS.n2568 VSS.n431 18.4216
R1245 VSS.n2569 VSS.n2568 18.4216
R1246 VSS.n2584 VSS.n421 18.4216
R1247 VSS.n2589 VSS.n421 18.4216
R1248 VSS.n2589 VSS.n419 18.4216
R1249 VSS.n2593 VSS.n419 18.4216
R1250 VSS.n2593 VSS.n416 18.4216
R1251 VSS.n2598 VSS.n416 18.4216
R1252 VSS.n2598 VSS.n414 18.4216
R1253 VSS.n2603 VSS.n414 18.4216
R1254 VSS.n2603 VSS.n412 18.4216
R1255 VSS.n2607 VSS.n412 18.4216
R1256 VSS.n2607 VSS.n409 18.4216
R1257 VSS.n2611 VSS.n409 18.4216
R1258 VSS.n2611 VSS.n407 18.4216
R1259 VSS.n2615 VSS.n407 18.4216
R1260 VSS.n2615 VSS.n405 18.4216
R1261 VSS.n2619 VSS.n405 18.4216
R1262 VSS.n2619 VSS.n402 18.4216
R1263 VSS.n2653 VSS.n402 18.4216
R1264 VSS.n2659 VSS.n399 18.4216
R1265 VSS.n2659 VSS.n397 18.4216
R1266 VSS.n2663 VSS.n397 18.4216
R1267 VSS.n2664 VSS.n2663 18.4216
R1268 VSS.n2664 VSS.n393 18.4216
R1269 VSS.n2696 VSS.n393 18.4216
R1270 VSS.n2696 VSS.n395 18.4216
R1271 VSS.n2692 VSS.n395 18.4216
R1272 VSS.n2692 VSS.n2668 18.4216
R1273 VSS.n2688 VSS.n2668 18.4216
R1274 VSS.n2688 VSS.n2670 18.4216
R1275 VSS.n2684 VSS.n2670 18.4216
R1276 VSS.n2684 VSS.n2672 18.4216
R1277 VSS.n2680 VSS.n2672 18.4216
R1278 VSS.n2680 VSS.n2674 18.4216
R1279 VSS.n2676 VSS.n2674 18.4216
R1280 VSS.n2676 VSS.n122 18.4216
R1281 VSS.n3240 VSS.n122 18.4216
R1282 VSS.n738 VSS.n736 18.4216
R1283 VSS.n754 VSS.n731 18.4216
R1284 VSS.n754 VSS.n732 18.4216
R1285 VSS.n750 VSS.n749 18.4216
R1286 VSS.n746 VSS.n745 18.4216
R1287 VSS.n742 VSS.n727 18.4216
R1288 VSS.n758 VSS.n757 18.4216
R1289 VSS.n762 VSS.n761 18.4216
R1290 VSS.n3403 VSS.n22 18.4216
R1291 VSS.n3399 VSS.n22 18.4216
R1292 VSS.n3399 VSS.n25 18.4216
R1293 VSS.n3395 VSS.n25 18.4216
R1294 VSS.n3395 VSS.n27 18.4216
R1295 VSS.n3391 VSS.n27 18.4216
R1296 VSS.n3391 VSS.n29 18.4216
R1297 VSS.n3387 VSS.n29 18.4216
R1298 VSS.n3387 VSS.n31 18.4216
R1299 VSS.n3383 VSS.n31 18.4216
R1300 VSS.n3383 VSS.n33 18.4216
R1301 VSS.n3379 VSS.n33 18.4216
R1302 VSS.n3379 VSS.n35 18.4216
R1303 VSS.n3375 VSS.n35 18.4216
R1304 VSS.n3375 VSS.n37 18.4216
R1305 VSS.n3371 VSS.n37 18.4216
R1306 VSS.n3371 VSS.n39 18.4216
R1307 VSS.n3367 VSS.n39 18.4216
R1308 VSS.n3363 VSS.n44 18.4216
R1309 VSS.n3359 VSS.n44 18.4216
R1310 VSS.n3359 VSS.n47 18.4216
R1311 VSS.n3355 VSS.n47 18.4216
R1312 VSS.n3355 VSS.n49 18.4216
R1313 VSS.n3351 VSS.n49 18.4216
R1314 VSS.n3351 VSS.n51 18.4216
R1315 VSS.n3347 VSS.n51 18.4216
R1316 VSS.n3347 VSS.n53 18.4216
R1317 VSS.n3343 VSS.n53 18.4216
R1318 VSS.n3343 VSS.n55 18.4216
R1319 VSS.n3339 VSS.n55 18.4216
R1320 VSS.n3339 VSS.n57 18.4216
R1321 VSS.n3335 VSS.n57 18.4216
R1322 VSS.n3335 VSS.n59 18.4216
R1323 VSS.n3331 VSS.n59 18.4216
R1324 VSS.n3331 VSS.n61 18.4216
R1325 VSS.n3327 VSS.n61 18.4216
R1326 VSS.n3323 VSS.n66 18.4216
R1327 VSS.n3319 VSS.n66 18.4216
R1328 VSS.n3319 VSS.n69 18.4216
R1329 VSS.n3315 VSS.n69 18.4216
R1330 VSS.n3315 VSS.n71 18.4216
R1331 VSS.n3311 VSS.n71 18.4216
R1332 VSS.n3311 VSS.n73 18.4216
R1333 VSS.n3307 VSS.n73 18.4216
R1334 VSS.n3307 VSS.n75 18.4216
R1335 VSS.n3303 VSS.n75 18.4216
R1336 VSS.n3303 VSS.n77 18.4216
R1337 VSS.n3299 VSS.n77 18.4216
R1338 VSS.n3299 VSS.n79 18.4216
R1339 VSS.n3295 VSS.n79 18.4216
R1340 VSS.n3295 VSS.n81 18.4216
R1341 VSS.n3291 VSS.n81 18.4216
R1342 VSS.n3291 VSS.n83 18.4216
R1343 VSS.n3287 VSS.n83 18.4216
R1344 VSS.n3283 VSS.n88 18.4216
R1345 VSS.n3279 VSS.n88 18.4216
R1346 VSS.n3279 VSS.n91 18.4216
R1347 VSS.n3275 VSS.n91 18.4216
R1348 VSS.n3275 VSS.n93 18.4216
R1349 VSS.n3271 VSS.n93 18.4216
R1350 VSS.n3271 VSS.n94 18.4216
R1351 VSS.n3267 VSS.n94 18.4216
R1352 VSS.n3267 VSS.n96 18.4216
R1353 VSS.n204 VSS.n96 18.4216
R1354 VSS.n207 VSS.n204 18.4216
R1355 VSS.n207 VSS.n203 18.4216
R1356 VSS.n211 VSS.n203 18.4216
R1357 VSS.n211 VSS.n201 18.4216
R1358 VSS.n216 VSS.n201 18.4216
R1359 VSS.n216 VSS.n199 18.4216
R1360 VSS.n220 VSS.n199 18.4216
R1361 VSS.n221 VSS.n220 18.4216
R1362 VSS.n2818 VSS.n197 18.4216
R1363 VSS.n2814 VSS.n197 18.4216
R1364 VSS.n2814 VSS.n225 18.4216
R1365 VSS.n2810 VSS.n225 18.4216
R1366 VSS.n2810 VSS.n227 18.4216
R1367 VSS.n2806 VSS.n227 18.4216
R1368 VSS.n2806 VSS.n229 18.4216
R1369 VSS.n2802 VSS.n229 18.4216
R1370 VSS.n2802 VSS.n231 18.4216
R1371 VSS.n2798 VSS.n231 18.4216
R1372 VSS.n2798 VSS.n233 18.4216
R1373 VSS.n2794 VSS.n233 18.4216
R1374 VSS.n2794 VSS.n235 18.4216
R1375 VSS.n2790 VSS.n235 18.4216
R1376 VSS.n2790 VSS.n237 18.4216
R1377 VSS.n2786 VSS.n237 18.4216
R1378 VSS.n2786 VSS.n238 18.4216
R1379 VSS.n2782 VSS.n238 18.4216
R1380 VSS.n2778 VSS.n2774 18.4216
R1381 VSS.n2774 VSS.n163 18.4216
R1382 VSS.n3118 VSS.n163 18.4216
R1383 VSS.n3120 VSS.n3118 18.4216
R1384 VSS.n3124 VSS.n161 18.4216
R1385 VSS.n3125 VSS.n3124 18.4216
R1386 VSS.n3127 VSS.n159 18.4216
R1387 VSS.n3131 VSS.n159 18.4216
R1388 VSS.n3134 VSS.n3133 18.4216
R1389 VSS.n3136 VSS.n3134 18.4216
R1390 VSS.n3140 VSS.n156 18.4216
R1391 VSS.n3143 VSS.n3142 18.4216
R1392 VSS.n3153 VSS.n3151 18.4216
R1393 VSS.n3157 VSS.n150 18.4216
R1394 VSS.n3161 VSS.n3159 18.4216
R1395 VSS.n3165 VSS.n148 18.4216
R1396 VSS.n3169 VSS.n3167 18.4216
R1397 VSS.n3173 VSS.n146 18.4216
R1398 VSS.n3177 VSS.n3175 18.4216
R1399 VSS.n3181 VSS.n144 18.4216
R1400 VSS.n3184 VSS.n3183 18.4216
R1401 VSS.n315 VSS.n314 18.4216
R1402 VSS.n318 VSS.n315 18.4216
R1403 VSS.n318 VSS.n311 18.4216
R1404 VSS.n322 VSS.n311 18.4216
R1405 VSS.n322 VSS.n309 18.4216
R1406 VSS.n327 VSS.n308 18.4216
R1407 VSS.n333 VSS.n308 18.4216
R1408 VSS.n335 VSS.n333 18.4216
R1409 VSS.n339 VSS.n306 18.4216
R1410 VSS.n343 VSS.n341 18.4216
R1411 VSS.n347 VSS.n304 18.4216
R1412 VSS.n364 VSS.n363 18.4216
R1413 VSS.n361 VSS.n352 18.4216
R1414 VSS.n357 VSS.n356 18.4216
R1415 VSS.n2706 VSS.n288 18.4216
R1416 VSS.n2706 VSS.n289 18.4216
R1417 VSS.n2702 VSS.n289 18.4216
R1418 VSS.n2702 VSS.n292 18.4216
R1419 VSS.n2630 VSS.n292 18.4216
R1420 VSS.n2631 VSS.n2630 18.4216
R1421 VSS.n2632 VSS.n2631 18.4216
R1422 VSS.n2639 VSS.n2638 18.4216
R1423 VSS.n2643 VSS.n2642 18.4216
R1424 VSS.n2647 VSS.n2626 18.4216
R1425 VSS.n1783 VSS.n918 18.4216
R1426 VSS.n1779 VSS.n918 18.4216
R1427 VSS.n1779 VSS.n1778 18.4216
R1428 VSS.n1778 VSS.n1734 18.4216
R1429 VSS.n1774 VSS.n1734 18.4216
R1430 VSS.n1774 VSS.n1736 18.4216
R1431 VSS.n1770 VSS.n1736 18.4216
R1432 VSS.n1770 VSS.n1739 18.4216
R1433 VSS.n1766 VSS.n1739 18.4216
R1434 VSS.n1766 VSS.n1741 18.4216
R1435 VSS.n1762 VSS.n1741 18.4216
R1436 VSS.n1762 VSS.n1743 18.4216
R1437 VSS.n1758 VSS.n1743 18.4216
R1438 VSS.n1758 VSS.n1745 18.4216
R1439 VSS.n1754 VSS.n1745 18.4216
R1440 VSS.n1754 VSS.n1747 18.4216
R1441 VSS.n1750 VSS.n1747 18.4216
R1442 VSS.n1750 VSS.n834 18.4216
R1443 VSS.n886 VSS.n835 18.4216
R1444 VSS.n882 VSS.n835 18.4216
R1445 VSS.n882 VSS.n838 18.4216
R1446 VSS.n878 VSS.n838 18.4216
R1447 VSS.n878 VSS.n841 18.4216
R1448 VSS.n874 VSS.n841 18.4216
R1449 VSS.n874 VSS.n843 18.4216
R1450 VSS.n870 VSS.n843 18.4216
R1451 VSS.n870 VSS.n845 18.4216
R1452 VSS.n866 VSS.n845 18.4216
R1453 VSS.n866 VSS.n847 18.4216
R1454 VSS.n862 VSS.n847 18.4216
R1455 VSS.n862 VSS.n849 18.4216
R1456 VSS.n858 VSS.n849 18.4216
R1457 VSS.n858 VSS.n851 18.4216
R1458 VSS.n854 VSS.n851 18.4216
R1459 VSS.n854 VSS.n716 18.4216
R1460 VSS.n2063 VSS.n716 18.4216
R1461 VSS.n2068 VSS.n2065 18.4216
R1462 VSS.n2068 VSS.n712 18.4216
R1463 VSS.n2072 VSS.n712 18.4216
R1464 VSS.n2072 VSS.n710 18.4216
R1465 VSS.n2076 VSS.n710 18.4216
R1466 VSS.n2076 VSS.n708 18.4216
R1467 VSS.n2080 VSS.n708 18.4216
R1468 VSS.n2080 VSS.n706 18.4216
R1469 VSS.n2084 VSS.n706 18.4216
R1470 VSS.n2084 VSS.n704 18.4216
R1471 VSS.n2088 VSS.n704 18.4216
R1472 VSS.n2088 VSS.n702 18.4216
R1473 VSS.n2092 VSS.n702 18.4216
R1474 VSS.n2092 VSS.n700 18.4216
R1475 VSS.n2097 VSS.n700 18.4216
R1476 VSS.n2097 VSS.n697 18.4216
R1477 VSS.n2101 VSS.n697 18.4216
R1478 VSS.n2102 VSS.n2101 18.4216
R1479 VSS.n2153 VSS.n2104 18.4216
R1480 VSS.n2149 VSS.n2104 18.4216
R1481 VSS.n2149 VSS.n2106 18.4216
R1482 VSS.n2145 VSS.n2106 18.4216
R1483 VSS.n2145 VSS.n2108 18.4216
R1484 VSS.n2141 VSS.n2108 18.4216
R1485 VSS.n2141 VSS.n2110 18.4216
R1486 VSS.n2137 VSS.n2110 18.4216
R1487 VSS.n2137 VSS.n2112 18.4216
R1488 VSS.n2133 VSS.n2112 18.4216
R1489 VSS.n2133 VSS.n2114 18.4216
R1490 VSS.n2129 VSS.n2114 18.4216
R1491 VSS.n2129 VSS.n2116 18.4216
R1492 VSS.n2125 VSS.n2116 18.4216
R1493 VSS.n2125 VSS.n2118 18.4216
R1494 VSS.n2121 VSS.n2118 18.4216
R1495 VSS.n2121 VSS.n537 18.4216
R1496 VSS.n2340 VSS.n537 18.4216
R1497 VSS.n2345 VSS.n2342 18.4216
R1498 VSS.n2345 VSS.n533 18.4216
R1499 VSS.n2349 VSS.n533 18.4216
R1500 VSS.n2349 VSS.n531 18.4216
R1501 VSS.n2353 VSS.n531 18.4216
R1502 VSS.n2353 VSS.n529 18.4216
R1503 VSS.n2357 VSS.n529 18.4216
R1504 VSS.n2357 VSS.n527 18.4216
R1505 VSS.n2361 VSS.n527 18.4216
R1506 VSS.n2361 VSS.n525 18.4216
R1507 VSS.n2365 VSS.n525 18.4216
R1508 VSS.n2365 VSS.n523 18.4216
R1509 VSS.n2369 VSS.n523 18.4216
R1510 VSS.n2369 VSS.n521 18.4216
R1511 VSS.n2374 VSS.n521 18.4216
R1512 VSS.n2374 VSS.n519 18.4216
R1513 VSS.n2378 VSS.n519 18.4216
R1514 VSS.n2379 VSS.n2378 18.4216
R1515 VSS.n2483 VSS.n2482 18.4216
R1516 VSS.n2482 VSS.n2382 18.4216
R1517 VSS.n2478 VSS.n2382 18.4216
R1518 VSS.n2478 VSS.n2384 18.4216
R1519 VSS.n2474 VSS.n2384 18.4216
R1520 VSS.n2474 VSS.n2387 18.4216
R1521 VSS.n2470 VSS.n2387 18.4216
R1522 VSS.n2470 VSS.n2389 18.4216
R1523 VSS.n2466 VSS.n2389 18.4216
R1524 VSS.n2466 VSS.n2391 18.4216
R1525 VSS.n2462 VSS.n2391 18.4216
R1526 VSS.n2462 VSS.n2393 18.4216
R1527 VSS.n2458 VSS.n2393 18.4216
R1528 VSS.n2458 VSS.n2395 18.4216
R1529 VSS.n2454 VSS.n2395 18.4216
R1530 VSS.n2454 VSS.n2397 18.4216
R1531 VSS.n2450 VSS.n2397 18.4216
R1532 VSS.n2450 VSS.n2398 18.4216
R1533 VSS.n2744 VSS.n264 18.4216
R1534 VSS.n2740 VSS.n264 18.4216
R1535 VSS.n2740 VSS.n266 18.4216
R1536 VSS.n2736 VSS.n266 18.4216
R1537 VSS.n2734 VSS.n2733 18.4216
R1538 VSS.n2731 VSS.n270 18.4216
R1539 VSS.n2727 VSS.n270 18.4216
R1540 VSS.n2727 VSS.n272 18.4216
R1541 VSS.n2723 VSS.n272 18.4216
R1542 VSS.n2723 VSS.n279 18.4216
R1543 VSS.n2719 VSS.n279 18.4216
R1544 VSS.n2719 VSS.n281 18.4216
R1545 VSS.n2715 VSS.n281 18.4216
R1546 VSS.n2715 VSS.n283 18.4216
R1547 VSS.n2711 VSS.n283 18.4216
R1548 VSS.n2711 VSS.n285 18.4216
R1549 VSS.n371 VSS.n301 18.4216
R1550 VSS.n371 VSS.n299 18.4216
R1551 VSS.n375 VSS.n299 18.4216
R1552 VSS.n375 VSS.n296 18.4216
R1553 VSS.n389 VSS.n296 18.4216
R1554 VSS.n389 VSS.n297 18.4216
R1555 VSS.n385 VSS.n297 18.4216
R1556 VSS.n385 VSS.n379 18.4216
R1557 VSS.n381 VSS.n379 18.4216
R1558 VSS.n381 VSS.n133 18.4216
R1559 VSS.n3220 VSS.n133 18.4216
R1560 VSS.n3220 VSS.n134 18.4216
R1561 VSS.n3216 VSS.n134 18.4216
R1562 VSS.n3214 VSS.n3213 18.4216
R1563 VSS.n3211 VSS.n138 18.4216
R1564 VSS.n1849 VSS.n1844 18.4216
R1565 VSS.n1865 VSS.n1841 18.4216
R1566 VSS.n1865 VSS.n1842 18.4216
R1567 VSS.n1861 VSS.n1860 18.4216
R1568 VSS.n1857 VSS.n1856 18.4216
R1569 VSS.n1853 VSS.n888 18.4216
R1570 VSS.n1869 VSS.n1868 18.4216
R1571 VSS.n1873 VSS.n1872 18.4216
R1572 VSS.n1887 VSS.n1886 17.4841
R1573 VSS.n2061 VSS.n2060 17.4841
R1574 VSS.n2164 VSS.n2163 17.4841
R1575 VSS.n2338 VSS.n2337 17.4841
R1576 VSS.n2489 VSS.n191 17.4841
R1577 VSS.n1169 VSS.n1016 16.9479
R1578 VSS.n1120 VSS.n1019 16.9479
R1579 VSS.n1713 VSS.t22 16.926
R1580 VSS.n1121 VSS.n1112 16.5247
R1581 VSS.n2822 VSS.n188 16.1749
R1582 VSS.t14 VSS.n2796 16.1749
R1583 VSS.t27 VSS.t54 15.6666
R1584 VSS.n3204 VSS.n141 15.0319
R1585 VSS.n1223 VSS.n992 14.5036
R1586 VSS.n1184 VSS.n1183 13.8958
R1587 VSS.n1712 VSS.t267 13.8486
R1588 VSS.n3256 VSS.n109 13.706
R1589 VSS.n1561 VSS.n1560 13.676
R1590 VSS.n1233 VSS.n1232 13.5743
R1591 VSS.n3262 VSS.n103 13.0685
R1592 VSS.n97 VSS.t0 12.9931
R1593 VSS.n1877 VSS.n886 12.5268
R1594 VSS.n2065 VSS.n2064 12.5268
R1595 VSS.n2153 VSS.n2103 12.5268
R1596 VSS.n2342 VSS.n2341 12.5268
R1597 VSS.n2483 VSS.n478 12.5268
R1598 VSS.n2744 VSS.n260 12.5268
R1599 VSS.n350 VSS.n301 12.5268
R1600 VSS.n3428 VSS.n3427 12.4628
R1601 VSS.n2822 VSS.n2821 12.4628
R1602 VSS.n1633 VSS.t262 12.4059
R1603 VSS.n1944 VSS.t190 12.4059
R1604 VSS.n1978 VSS.t220 12.4059
R1605 VSS.n2221 VSS.t194 12.4059
R1606 VSS.n2255 VSS.t192 12.4059
R1607 VSS.n440 VSS.t260 12.4059
R1608 VSS.n410 VSS.t122 12.3005
R1609 VSS.n954 VSS.n942 12.033
R1610 VSS.n1691 VSS.n1685 12.033
R1611 VSS.n1691 VSS.n1684 12.033
R1612 VSS.n3258 VSS.t217 11.9233
R1613 VSS.n2699 VSS.n2698 11.6366
R1614 VSS.n129 VSS.n125 11.4244
R1615 VSS.n1929 VSS.n807 11.4216
R1616 VSS.n2021 VSS.n787 11.4216
R1617 VSS.n2206 VSS.n628 11.4216
R1618 VSS.n2298 VSS.n608 11.4216
R1619 VSS.n452 VSS.n448 11.4216
R1620 VSS.n2584 VSS.n423 11.4216
R1621 VSS.n403 VSS.n399 11.4216
R1622 VSS.n3363 VSS.n41 11.4216
R1623 VSS.n3323 VSS.n63 11.4216
R1624 VSS.n3283 VSS.n85 11.4216
R1625 VSS.n2818 VSS.n196 11.4216
R1626 VSS.n2778 VSS.n240 11.4216
R1627 VSS.n3149 VSS.n152 11.4216
R1628 VSS.n3237 VSS.n119 11.3366
R1629 VSS.n104 VSS.t44 11.1395
R1630 VSS.n956 VSS.t34 11.0292
R1631 VSS.n1690 VSS.t252 11.0292
R1632 VSS.n1690 VSS.t114 11.0292
R1633 VSS.n1075 VSS.t53 11.0225
R1634 VSS.n141 VSS.n108 10.6137
R1635 VSS.t13 VSS.n3265 10.6067
R1636 VSS.n1718 VSS.t230 10.5091
R1637 VSS.n1205 VSS.n1076 10.4005
R1638 VSS.n1204 VSS.n1203 10.4005
R1639 VSS.n1202 VSS.n1201 10.4005
R1640 VSS.n1084 VSS.n1083 10.4005
R1641 VSS.t52 VSS.n1074 10.4005
R1642 VSS.n1085 VSS.t104 10.4005
R1643 VSS.t59 VSS.n1200 10.4005
R1644 VSS.n1199 VSS.t45 10.4005
R1645 VSS.n1234 VSS.n1233 10.4005
R1646 VSS.n1562 VSS.n1561 10.4005
R1647 VSS.n3116 VSS.n173 10.4005
R1648 VSS.n3116 VSS.n172 10.4005
R1649 VSS.n3116 VSS.n174 10.4005
R1650 VSS.n3116 VSS.n171 10.4005
R1651 VSS.n3116 VSS.n175 10.4005
R1652 VSS.n3116 VSS.n170 10.4005
R1653 VSS.n3116 VSS.n176 10.4005
R1654 VSS.n3116 VSS.n169 10.4005
R1655 VSS.n3116 VSS.n177 10.4005
R1656 VSS.n3116 VSS.n168 10.4005
R1657 VSS.n3116 VSS.n178 10.4005
R1658 VSS.n3116 VSS.n167 10.4005
R1659 VSS.n3116 VSS.n179 10.4005
R1660 VSS.n3116 VSS.n166 10.4005
R1661 VSS.n3116 VSS.n180 10.4005
R1662 VSS.n3116 VSS.n165 10.4005
R1663 VSS.n3116 VSS.n3115 10.4005
R1664 VSS.n931 VSS.t92 10.2792
R1665 VSS.n1704 VSS.t94 10.2607
R1666 VSS.n1719 VSS.t176 10.0514
R1667 VSS.n1721 VSS.t180 10.0514
R1668 VSS.t129 VSS.t269 9.96983
R1669 VSS.n1116 VSS.n1115 9.94787
R1670 VSS.n1182 VSS.n1181 9.94787
R1671 VSS.n1925 VSS.n807 9.94787
R1672 VSS.n1967 VSS.n787 9.94787
R1673 VSS.n2202 VSS.n628 9.94787
R1674 VSS.n2244 VSS.n608 9.94787
R1675 VSS.n2529 VSS.n452 9.94787
R1676 VSS.n2569 VSS.n423 9.94787
R1677 VSS.n2653 VSS.n403 9.94787
R1678 VSS.n3367 VSS.n41 9.94787
R1679 VSS.n3327 VSS.n63 9.94787
R1680 VSS.n3287 VSS.n85 9.94787
R1681 VSS.n221 VSS.n196 9.94787
R1682 VSS.n2782 VSS.n240 9.94787
R1683 VSS.n3145 VSS.n152 9.94787
R1684 VSS.n972 VSS.t166 9.93604
R1685 VSS.n976 VSS.t57 9.93604
R1686 VSS.n979 VSS.t119 9.93604
R1687 VSS.n989 VSS.t112 9.93604
R1688 VSS.n946 VSS.t139 9.93604
R1689 VSS.n951 VSS.t143 9.93604
R1690 VSS.n952 VSS.t78 9.93604
R1691 VSS.n960 VSS.t64 9.93604
R1692 VSS.n960 VSS.t63 9.93604
R1693 VSS.n1674 VSS.n933 9.73801
R1694 VSS.n1887 VSS.n23 9.71359
R1695 VSS.n2060 VSS.n45 9.71359
R1696 VSS.n2164 VSS.n67 9.71359
R1697 VSS.n2337 VSS.n89 9.71359
R1698 VSS.n2820 VSS.n191 9.71359
R1699 VSS.n3225 VSS.n129 9.188
R1700 VSS.n1722 VSS.t172 9.15882
R1701 VSS.n3195 VSS.t202 9.05408
R1702 VSS.n1783 VSS.n917 9.02682
R1703 VSS.t45 VSS.n1084 9.01367
R1704 VSS.n3259 VSS.n3258 8.92063
R1705 VSS.n1877 VSS.n834 8.84261
R1706 VSS.n2064 VSS.n2063 8.84261
R1707 VSS.n2103 VSS.n2102 8.84261
R1708 VSS.n2341 VSS.n2340 8.84261
R1709 VSS.n2379 VSS.n478 8.84261
R1710 VSS.n2398 VSS.n260 8.84261
R1711 VSS.n350 VSS.n285 8.84261
R1712 VSS.n2824 VSS.n2823 8.77991
R1713 VSS.n966 VSS.t145 8.51132
R1714 VSS.n1215 VSS.t283 8.51132
R1715 VSS.n1216 VSS.t273 8.51132
R1716 VSS.n1217 VSS.t124 8.51132
R1717 VSS.n1218 VSS.t55 8.51132
R1718 VSS.n1220 VSS.t281 8.51132
R1719 VSS.n1221 VSS.t51 8.51132
R1720 VSS.n1214 VSS.t155 8.51132
R1721 VSS.n1213 VSS.t42 8.51132
R1722 VSS.n988 VSS.t159 8.51132
R1723 VSS.n986 VSS.t61 8.51132
R1724 VSS.n984 VSS.t12 8.51132
R1725 VSS.n983 VSS.t66 8.51132
R1726 VSS.n981 VSS.t18 8.51132
R1727 VSS.n978 VSS.t293 8.51132
R1728 VSS.n939 VSS.t16 8.51132
R1729 VSS.n1696 VSS.t211 8.51132
R1730 VSS.n1688 VSS.t297 8.51132
R1731 VSS.n1688 VSS.t148 8.51132
R1732 VSS.n1697 VSS.t218 8.51132
R1733 VSS.n975 VSS.t76 8.48197
R1734 VSS.n948 VSS.t49 8.46241
R1735 VSS.n1693 VSS.t72 8.46241
R1736 VSS.n1693 VSS.t258 8.46241
R1737 VSS.n974 VSS.t256 8.4135
R1738 VSS.n982 VSS.t289 8.4135
R1739 VSS.n985 VSS.t116 8.4135
R1740 VSS.n987 VSS.t4 8.4135
R1741 VSS.n949 VSS.t82 8.4135
R1742 VSS.n955 VSS.t266 8.4135
R1743 VSS.n957 VSS.t80 8.4135
R1744 VSS.n959 VSS.t285 8.4135
R1745 VSS.n942 VSS.t251 8.4005
R1746 VSS.n942 VSS.t2 8.4005
R1747 VSS.n1685 VSS.t149 8.4005
R1748 VSS.n1685 VSS.t68 8.4005
R1749 VSS.n1684 VSS.t6 8.4005
R1750 VSS.n1684 VSS.t301 8.4005
R1751 VSS.n3204 VSS.n3203 8.28675
R1752 VSS.n3403 VSS.n21 8.14755
R1753 VSS.n944 VSS.t47 8.0855
R1754 VSS.n1683 VSS.t70 8.0855
R1755 VSS.n1682 VSS.t257 8.0855
R1756 VSS.n1921 VSS.n807 7.92155
R1757 VSS.n2025 VSS.n787 7.92155
R1758 VSS.n2198 VSS.n628 7.92155
R1759 VSS.n2302 VSS.n608 7.92155
R1760 VSS.n455 VSS.n452 7.92155
R1761 VSS.n2580 VSS.n423 7.92155
R1762 VSS.n2648 VSS.n403 7.92155
R1763 VSS.n1878 VSS.n1877 7.82945
R1764 VSS.n2064 VSS.n714 7.82945
R1765 VSS.n2103 VSS.n653 7.82945
R1766 VSS.n2341 VSS.n536 7.82945
R1767 VSS.n516 VSS.n478 7.82945
R1768 VSS.n2403 VSS.n260 7.82945
R1769 VSS.n366 VSS.n350 7.82945
R1770 VSS.n1179 VSS.n1109 7.74316
R1771 VSS.n1495 VSS.n1016 7.36892
R1772 VSS.n1493 VSS.n1019 7.36892
R1773 VSS.n1106 VSS.t38 7.13593
R1774 VSS.n1180 VSS.t36 7.13593
R1775 VSS.n3203 VSS.n128 7.1055
R1776 VSS.n1710 VSS.n935 6.94217
R1777 VSS.n241 VSS.n194 6.62937
R1778 VSS.n125 VSS.n123 6.62351
R1779 VSS.n950 VSS.n944 6.54898
R1780 VSS.n1692 VSS.n1682 6.54898
R1781 VSS.n1692 VSS.n1683 6.54898
R1782 VSS.n958 VSS.n941 6.46859
R1783 VSS.n1689 VSS.n1686 6.46859
R1784 VSS.n1689 VSS.n1687 6.46859
R1785 VSS.n1717 VSS.n930 6.46462
R1786 VSS.n1703 VSS.n1698 6.45138
R1787 VSS.n1702 VSS.n1699 6.45138
R1788 VSS.n1701 VSS.n1700 6.45138
R1789 VSS.n1720 VSS.n929 6.45138
R1790 VSS.n245 VSS.n240 6.44787
R1791 VSS.n484 VSS.n196 6.44787
R1792 VSS.n555 VSS.n85 6.44787
R1793 VSS.n663 VSS.n63 6.44787
R1794 VSS.n734 VSS.n41 6.44787
R1795 VSS.n3184 VSS.n102 6.44787
R1796 VSS.n314 VSS.n152 6.44787
R1797 VSS.n1845 VSS.n21 6.44787
R1798 VSS.n1211 VSS.t128 6.3005
R1799 VSS.n1205 VSS.t52 6.00928
R1800 VSS.n916 VSS.n889 5.82835
R1801 VSS.n1211 VSS.t305 5.6196
R1802 VSS.n1590 VSS.n889 5.5943
R1803 VSS.n3261 VSS.n3260 5.39487
R1804 VSS.n3207 VSS.n3206 5.34261
R1805 VSS.n1555 VSS.n1554 5.32359
R1806 VSS.n1209 VSS.n937 5.32359
R1807 VSS.n977 VSS.n968 5.32359
R1808 VSS.n973 VSS.n969 5.32359
R1809 VSS.n971 VSS.n970 5.32359
R1810 VSS.n938 VSS.n934 5.32359
R1811 VSS.n947 VSS.n945 5.32359
R1812 VSS.n1695 VSS.n940 5.32359
R1813 VSS.n990 VSS.n963 5.32226
R1814 VSS.n980 VSS.n967 5.32226
R1815 VSS.n953 VSS.n943 5.32226
R1816 VSS.n1694 VSS.n1681 5.32226
R1817 VSS.n1723 VSS.n928 5.32226
R1818 VSS.n2698 VSS.n393 5.23035
R1819 VSS.n1196 VSS.n1086 5.2014
R1820 VSS.n1915 VSS.n814 5.2005
R1821 VSS.n1915 VSS.n1914 5.2005
R1822 VSS.n1909 VSS.n815 5.2005
R1823 VSS.n1913 VSS.n815 5.2005
R1824 VSS.n1911 VSS.n1910 5.2005
R1825 VSS.n1912 VSS.n1911 5.2005
R1826 VSS.n1908 VSS.n817 5.2005
R1827 VSS.n817 VSS.n816 5.2005
R1828 VSS.n1907 VSS.n1906 5.2005
R1829 VSS.n1906 VSS.n1905 5.2005
R1830 VSS.n819 VSS.n818 5.2005
R1831 VSS.n1904 VSS.n819 5.2005
R1832 VSS.n1902 VSS.n1901 5.2005
R1833 VSS.n1903 VSS.n1902 5.2005
R1834 VSS.n1900 VSS.n821 5.2005
R1835 VSS.n821 VSS.n820 5.2005
R1836 VSS.n1899 VSS.n1898 5.2005
R1837 VSS.n1898 VSS.n1897 5.2005
R1838 VSS.n823 VSS.n822 5.2005
R1839 VSS.n1896 VSS.n823 5.2005
R1840 VSS.n1894 VSS.n1893 5.2005
R1841 VSS.n1895 VSS.n1894 5.2005
R1842 VSS.n1892 VSS.n825 5.2005
R1843 VSS.n825 VSS.n824 5.2005
R1844 VSS.n1891 VSS.n1890 5.2005
R1845 VSS.n1890 VSS.n1889 5.2005
R1846 VSS.n827 VSS.n826 5.2005
R1847 VSS.n1888 VSS.n827 5.2005
R1848 VSS.n2032 VSS.n783 5.2005
R1849 VSS.n783 VSS.n782 5.2005
R1850 VSS.n2034 VSS.n2033 5.2005
R1851 VSS.n2035 VSS.n2034 5.2005
R1852 VSS.n781 VSS.n780 5.2005
R1853 VSS.n2036 VSS.n781 5.2005
R1854 VSS.n2039 VSS.n2038 5.2005
R1855 VSS.n2038 VSS.n2037 5.2005
R1856 VSS.n2040 VSS.n779 5.2005
R1857 VSS.n779 VSS.n778 5.2005
R1858 VSS.n2042 VSS.n2041 5.2005
R1859 VSS.n2043 VSS.n2042 5.2005
R1860 VSS.n777 VSS.n776 5.2005
R1861 VSS.n2044 VSS.n777 5.2005
R1862 VSS.n2047 VSS.n2046 5.2005
R1863 VSS.n2046 VSS.n2045 5.2005
R1864 VSS.n2048 VSS.n775 5.2005
R1865 VSS.n775 VSS.n774 5.2005
R1866 VSS.n2050 VSS.n2049 5.2005
R1867 VSS.n2051 VSS.n2050 5.2005
R1868 VSS.n773 VSS.n772 5.2005
R1869 VSS.n2052 VSS.n773 5.2005
R1870 VSS.n2055 VSS.n2054 5.2005
R1871 VSS.n2054 VSS.n2053 5.2005
R1872 VSS.n2056 VSS.n725 5.2005
R1873 VSS.n725 VSS.n723 5.2005
R1874 VSS.n2058 VSS.n2057 5.2005
R1875 VSS.n2059 VSS.n2058 5.2005
R1876 VSS.n2192 VSS.n635 5.2005
R1877 VSS.n2192 VSS.n2191 5.2005
R1878 VSS.n2186 VSS.n636 5.2005
R1879 VSS.n2190 VSS.n636 5.2005
R1880 VSS.n2188 VSS.n2187 5.2005
R1881 VSS.n2189 VSS.n2188 5.2005
R1882 VSS.n2185 VSS.n638 5.2005
R1883 VSS.n638 VSS.n637 5.2005
R1884 VSS.n2184 VSS.n2183 5.2005
R1885 VSS.n2183 VSS.n2182 5.2005
R1886 VSS.n640 VSS.n639 5.2005
R1887 VSS.n2181 VSS.n640 5.2005
R1888 VSS.n2179 VSS.n2178 5.2005
R1889 VSS.n2180 VSS.n2179 5.2005
R1890 VSS.n2177 VSS.n642 5.2005
R1891 VSS.n642 VSS.n641 5.2005
R1892 VSS.n2176 VSS.n2175 5.2005
R1893 VSS.n2175 VSS.n2174 5.2005
R1894 VSS.n644 VSS.n643 5.2005
R1895 VSS.n2173 VSS.n644 5.2005
R1896 VSS.n2171 VSS.n2170 5.2005
R1897 VSS.n2172 VSS.n2171 5.2005
R1898 VSS.n2169 VSS.n646 5.2005
R1899 VSS.n646 VSS.n645 5.2005
R1900 VSS.n2168 VSS.n2167 5.2005
R1901 VSS.n2167 VSS.n2166 5.2005
R1902 VSS.n648 VSS.n647 5.2005
R1903 VSS.n2165 VSS.n648 5.2005
R1904 VSS.n2309 VSS.n604 5.2005
R1905 VSS.n604 VSS.n603 5.2005
R1906 VSS.n2311 VSS.n2310 5.2005
R1907 VSS.n2312 VSS.n2311 5.2005
R1908 VSS.n602 VSS.n601 5.2005
R1909 VSS.n2313 VSS.n602 5.2005
R1910 VSS.n2316 VSS.n2315 5.2005
R1911 VSS.n2315 VSS.n2314 5.2005
R1912 VSS.n2317 VSS.n600 5.2005
R1913 VSS.n600 VSS.n599 5.2005
R1914 VSS.n2319 VSS.n2318 5.2005
R1915 VSS.n2320 VSS.n2319 5.2005
R1916 VSS.n598 VSS.n597 5.2005
R1917 VSS.n2321 VSS.n598 5.2005
R1918 VSS.n2324 VSS.n2323 5.2005
R1919 VSS.n2323 VSS.n2322 5.2005
R1920 VSS.n2325 VSS.n596 5.2005
R1921 VSS.n596 VSS.n595 5.2005
R1922 VSS.n2327 VSS.n2326 5.2005
R1923 VSS.n2328 VSS.n2327 5.2005
R1924 VSS.n594 VSS.n593 5.2005
R1925 VSS.n2329 VSS.n594 5.2005
R1926 VSS.n2332 VSS.n2331 5.2005
R1927 VSS.n2331 VSS.n2330 5.2005
R1928 VSS.n2333 VSS.n546 5.2005
R1929 VSS.n546 VSS.n544 5.2005
R1930 VSS.n2335 VSS.n2334 5.2005
R1931 VSS.n2336 VSS.n2335 5.2005
R1932 VSS.n2524 VSS.n2523 5.2005
R1933 VSS.n2525 VSS.n2524 5.2005
R1934 VSS.n2517 VSS.n458 5.2005
R1935 VSS.n458 VSS.n457 5.2005
R1936 VSS.n2516 VSS.n2515 5.2005
R1937 VSS.n2515 VSS.n2514 5.2005
R1938 VSS.n461 VSS.n460 5.2005
R1939 VSS.n2513 VSS.n461 5.2005
R1940 VSS.n2511 VSS.n2510 5.2005
R1941 VSS.n2512 VSS.n2511 5.2005
R1942 VSS.n2509 VSS.n463 5.2005
R1943 VSS.n463 VSS.n462 5.2005
R1944 VSS.n2508 VSS.n2507 5.2005
R1945 VSS.n2507 VSS.n2506 5.2005
R1946 VSS.n465 VSS.n464 5.2005
R1947 VSS.n2505 VSS.n465 5.2005
R1948 VSS.n2503 VSS.n2502 5.2005
R1949 VSS.n2504 VSS.n2503 5.2005
R1950 VSS.n2501 VSS.n467 5.2005
R1951 VSS.n467 VSS.n466 5.2005
R1952 VSS.n2500 VSS.n2499 5.2005
R1953 VSS.n2499 VSS.n2498 5.2005
R1954 VSS.n469 VSS.n468 5.2005
R1955 VSS.n2497 VSS.n469 5.2005
R1956 VSS.n2495 VSS.n2494 5.2005
R1957 VSS.n2496 VSS.n2495 5.2005
R1958 VSS.n2493 VSS.n471 5.2005
R1959 VSS.n471 VSS.n470 5.2005
R1960 VSS.n1921 VSS.n808 5.2005
R1961 VSS.n1920 VSS.n1919 5.2005
R1962 VSS.n1918 VSS.n813 5.2005
R1963 VSS.n1917 VSS.n1916 5.2005
R1964 VSS.n2025 VSS.n2024 5.2005
R1965 VSS.n2027 VSS.n786 5.2005
R1966 VSS.n2028 VSS.n784 5.2005
R1967 VSS.n2031 VSS.n2030 5.2005
R1968 VSS.n2198 VSS.n629 5.2005
R1969 VSS.n2197 VSS.n2196 5.2005
R1970 VSS.n2195 VSS.n634 5.2005
R1971 VSS.n2194 VSS.n2193 5.2005
R1972 VSS.n2302 VSS.n2301 5.2005
R1973 VSS.n2304 VSS.n607 5.2005
R1974 VSS.n2305 VSS.n605 5.2005
R1975 VSS.n2308 VSS.n2307 5.2005
R1976 VSS.n455 VSS.n449 5.2005
R1977 VSS.n2519 VSS.n2518 5.2005
R1978 VSS.n2521 VSS.n2520 5.2005
R1979 VSS.n2522 VSS.n459 5.2005
R1980 VSS.n585 VSS.n535 5.2005
R1981 VSS.n584 VSS.n583 5.2005
R1982 VSS.n582 VSS.n581 5.2005
R1983 VSS.n580 VSS.n579 5.2005
R1984 VSS.n2487 VSS.n2486 5.2005
R1985 VSS.n513 VSS.n477 5.2005
R1986 VSS.n512 VSS.n511 5.2005
R1987 VSS.n510 VSS.n509 5.2005
R1988 VSS.n2748 VSS.n2747 5.2005
R1989 VSS.n2750 VSS.n257 5.2005
R1990 VSS.n2752 VSS.n2751 5.2005
R1991 VSS.n2753 VSS.n256 5.2005
R1992 VSS.n1884 VSS.n1883 5.2005
R1993 VSS.n1882 VSS.n832 5.2005
R1994 VSS.n1881 VSS.n1880 5.2005
R1995 VSS.n1879 VSS.n1878 5.2005
R1996 VSS.n771 VSS.n724 5.2005
R1997 VSS.n770 VSS.n769 5.2005
R1998 VSS.n768 VSS.n767 5.2005
R1999 VSS.n766 VSS.n714 5.2005
R2000 VSS.n2158 VSS.n2157 5.2005
R2001 VSS.n2159 VSS.n654 5.2005
R2002 VSS.n2161 VSS.n2160 5.2005
R2003 VSS.n2156 VSS.n653 5.2005
R2004 VSS.n592 VSS.n545 5.2005
R2005 VSS.n591 VSS.n590 5.2005
R2006 VSS.n589 VSS.n588 5.2005
R2007 VSS.n587 VSS.n536 5.2005
R2008 VSS.n2492 VSS.n2491 5.2005
R2009 VSS.n473 VSS.n472 5.2005
R2010 VSS.n515 VSS.n514 5.2005
R2011 VSS.n517 VSS.n516 5.2005
R2012 VSS.n696 VSS.n693 5.2005
R2013 VSS.n692 VSS.n691 5.2005
R2014 VSS.n690 VSS.n689 5.2005
R2015 VSS.n688 VSS.n687 5.2005
R2016 VSS.n686 VSS.n655 5.2005
R2017 VSS.n670 VSS.n656 5.2005
R2018 VSS.n672 VSS.n671 5.2005
R2019 VSS.n674 VSS.n673 5.2005
R2020 VSS.n676 VSS.n675 5.2005
R2021 VSS.n678 VSS.n677 5.2005
R2022 VSS.n680 VSS.n679 5.2005
R2023 VSS.n681 VSS.n661 5.2005
R2024 VSS.n683 VSS.n682 5.2005
R2025 VSS.n684 VSS.n683 5.2005
R2026 VSS.n578 VSS.n547 5.2005
R2027 VSS.n562 VSS.n548 5.2005
R2028 VSS.n564 VSS.n563 5.2005
R2029 VSS.n566 VSS.n565 5.2005
R2030 VSS.n568 VSS.n567 5.2005
R2031 VSS.n570 VSS.n569 5.2005
R2032 VSS.n572 VSS.n571 5.2005
R2033 VSS.n573 VSS.n553 5.2005
R2034 VSS.n575 VSS.n574 5.2005
R2035 VSS.n576 VSS.n575 5.2005
R2036 VSS.n508 VSS.n479 5.2005
R2037 VSS.n506 VSS.n505 5.2005
R2038 VSS.n504 VSS.n480 5.2005
R2039 VSS.n503 VSS.n502 5.2005
R2040 VSS.n500 VSS.n481 5.2005
R2041 VSS.n498 VSS.n497 5.2005
R2042 VSS.n496 VSS.n482 5.2005
R2043 VSS.n495 VSS.n494 5.2005
R2044 VSS.n492 VSS.n483 5.2005
R2045 VSS.n492 VSS.n193 5.2005
R2046 VSS.n2755 VSS.n2754 5.2005
R2047 VSS.n2757 VSS.n254 5.2005
R2048 VSS.n2759 VSS.n2758 5.2005
R2049 VSS.n2760 VSS.n253 5.2005
R2050 VSS.n2762 VSS.n2761 5.2005
R2051 VSS.n2764 VSS.n252 5.2005
R2052 VSS.n2765 VSS.n250 5.2005
R2053 VSS.n2768 VSS.n2767 5.2005
R2054 VSS.n2769 VSS.n244 5.2005
R2055 VSS.n251 VSS.n244 5.2005
R2056 VSS.n2581 VSS.n2580 5.2005
R2057 VSS.n2578 VSS.n425 5.2005
R2058 VSS.n2577 VSS.n2576 5.2005
R2059 VSS.n2575 VSS.n2574 5.2005
R2060 VSS.n2573 VSS.n427 5.2005
R2061 VSS.n2573 VSS.n2572 5.2005
R2062 VSS.n2421 VSS.n428 5.2005
R2063 VSS.n429 VSS.n428 5.2005
R2064 VSS.n2424 VSS.n2423 5.2005
R2065 VSS.n2423 VSS.n2422 5.2005
R2066 VSS.n2425 VSS.n2419 5.2005
R2067 VSS.n2419 VSS.n2418 5.2005
R2068 VSS.n2427 VSS.n2426 5.2005
R2069 VSS.n2428 VSS.n2427 5.2005
R2070 VSS.n2420 VSS.n2417 5.2005
R2071 VSS.n2429 VSS.n2417 5.2005
R2072 VSS.n2431 VSS.n2416 5.2005
R2073 VSS.n2431 VSS.n2430 5.2005
R2074 VSS.n2434 VSS.n2433 5.2005
R2075 VSS.n2433 VSS.n2432 5.2005
R2076 VSS.n2435 VSS.n2415 5.2005
R2077 VSS.n2415 VSS.n2414 5.2005
R2078 VSS.n2437 VSS.n2436 5.2005
R2079 VSS.n2438 VSS.n2437 5.2005
R2080 VSS.n2411 VSS.n2410 5.2005
R2081 VSS.n2439 VSS.n2411 5.2005
R2082 VSS.n2442 VSS.n2441 5.2005
R2083 VSS.n2441 VSS.n2440 5.2005
R2084 VSS.n2443 VSS.n2401 5.2005
R2085 VSS.n2401 VSS.n2399 5.2005
R2086 VSS.n2445 VSS.n2444 5.2005
R2087 VSS.n2446 VSS.n2445 5.2005
R2088 VSS.n2409 VSS.n2400 5.2005
R2089 VSS.n2408 VSS.n2407 5.2005
R2090 VSS.n2405 VSS.n2402 5.2005
R2091 VSS.n2403 VSS.n261 5.2005
R2092 VSS.n1674 VSS.n1673 5.2005
R2093 VSS.n1675 VSS.n1674 5.2005
R2094 VSS.n1672 VSS.n1572 5.2005
R2095 VSS.n1572 VSS.n1571 5.2005
R2096 VSS.n1671 VSS.n1670 5.2005
R2097 VSS.n1670 VSS.n1669 5.2005
R2098 VSS.n1575 VSS.n1574 5.2005
R2099 VSS.n1668 VSS.n1575 5.2005
R2100 VSS.n1666 VSS.n1665 5.2005
R2101 VSS.n1667 VSS.n1666 5.2005
R2102 VSS.n1664 VSS.n1628 5.2005
R2103 VSS.n1628 VSS.n1627 5.2005
R2104 VSS.n1663 VSS.n1662 5.2005
R2105 VSS.n1662 VSS.n1661 5.2005
R2106 VSS.n1630 VSS.n1629 5.2005
R2107 VSS.n1660 VSS.n1630 5.2005
R2108 VSS.n1658 VSS.n1657 5.2005
R2109 VSS.n1659 VSS.n1658 5.2005
R2110 VSS.n1655 VSS.n1632 5.2005
R2111 VSS.n1632 VSS.n1631 5.2005
R2112 VSS.n1654 VSS.n1653 5.2005
R2113 VSS.n1653 VSS.n1652 5.2005
R2114 VSS.n1635 VSS.n1634 5.2005
R2115 VSS.n1651 VSS.n1635 5.2005
R2116 VSS.n1649 VSS.n1648 5.2005
R2117 VSS.n1650 VSS.n1649 5.2005
R2118 VSS.n1647 VSS.n1637 5.2005
R2119 VSS.n1637 VSS.n1636 5.2005
R2120 VSS.n1646 VSS.n1645 5.2005
R2121 VSS.n1645 VSS.n1644 5.2005
R2122 VSS.n1639 VSS.n1638 5.2005
R2123 VSS.n1643 VSS.n1639 5.2005
R2124 VSS.n1641 VSS.n1640 5.2005
R2125 VSS.n1642 VSS.n1641 5.2005
R2126 VSS.n810 VSS.n809 5.2005
R2127 VSS.n811 VSS.n810 5.2005
R2128 VSS.n1926 VSS.n1925 5.2005
R2129 VSS.n1925 VSS.n1924 5.2005
R2130 VSS.n1929 VSS.n1928 5.2005
R2131 VSS.n1930 VSS.n1929 5.2005
R2132 VSS.n805 VSS.n804 5.2005
R2133 VSS.n1931 VSS.n805 5.2005
R2134 VSS.n1934 VSS.n1933 5.2005
R2135 VSS.n1933 VSS.n1932 5.2005
R2136 VSS.n1935 VSS.n803 5.2005
R2137 VSS.n803 VSS.n802 5.2005
R2138 VSS.n1937 VSS.n1936 5.2005
R2139 VSS.n1938 VSS.n1937 5.2005
R2140 VSS.n801 VSS.n800 5.2005
R2141 VSS.n1939 VSS.n801 5.2005
R2142 VSS.n1942 VSS.n1941 5.2005
R2143 VSS.n1941 VSS.n1940 5.2005
R2144 VSS.n1943 VSS.n799 5.2005
R2145 VSS.n799 VSS.n798 5.2005
R2146 VSS.n1947 VSS.n1946 5.2005
R2147 VSS.n1948 VSS.n1947 5.2005
R2148 VSS.n797 VSS.n796 5.2005
R2149 VSS.n1949 VSS.n797 5.2005
R2150 VSS.n1952 VSS.n1951 5.2005
R2151 VSS.n1951 VSS.n1950 5.2005
R2152 VSS.n1953 VSS.n795 5.2005
R2153 VSS.n795 VSS.n794 5.2005
R2154 VSS.n1955 VSS.n1954 5.2005
R2155 VSS.n1956 VSS.n1955 5.2005
R2156 VSS.n793 VSS.n792 5.2005
R2157 VSS.n1957 VSS.n793 5.2005
R2158 VSS.n1960 VSS.n1959 5.2005
R2159 VSS.n1959 VSS.n1958 5.2005
R2160 VSS.n1961 VSS.n791 5.2005
R2161 VSS.n791 VSS.n790 5.2005
R2162 VSS.n1963 VSS.n1962 5.2005
R2163 VSS.n1964 VSS.n1963 5.2005
R2164 VSS.n789 VSS.n788 5.2005
R2165 VSS.n1965 VSS.n789 5.2005
R2166 VSS.n1968 VSS.n1967 5.2005
R2167 VSS.n1967 VSS.n1966 5.2005
R2168 VSS.n2022 VSS.n2021 5.2005
R2169 VSS.n2021 VSS.n2020 5.2005
R2170 VSS.n1970 VSS.n1969 5.2005
R2171 VSS.n2019 VSS.n1970 5.2005
R2172 VSS.n2017 VSS.n2016 5.2005
R2173 VSS.n2018 VSS.n2017 5.2005
R2174 VSS.n2015 VSS.n1973 5.2005
R2175 VSS.n1973 VSS.n1972 5.2005
R2176 VSS.n2014 VSS.n2013 5.2005
R2177 VSS.n2013 VSS.n2012 5.2005
R2178 VSS.n1975 VSS.n1974 5.2005
R2179 VSS.n2011 VSS.n1975 5.2005
R2180 VSS.n2009 VSS.n2008 5.2005
R2181 VSS.n2010 VSS.n2009 5.2005
R2182 VSS.n2007 VSS.n1977 5.2005
R2183 VSS.n1977 VSS.n1976 5.2005
R2184 VSS.n2006 VSS.n2005 5.2005
R2185 VSS.n2005 VSS.n2004 5.2005
R2186 VSS.n1983 VSS.n1980 5.2005
R2187 VSS.n2003 VSS.n1980 5.2005
R2188 VSS.n2001 VSS.n2000 5.2005
R2189 VSS.n2002 VSS.n2001 5.2005
R2190 VSS.n1999 VSS.n1982 5.2005
R2191 VSS.n1982 VSS.n1981 5.2005
R2192 VSS.n1998 VSS.n1997 5.2005
R2193 VSS.n1997 VSS.n1996 5.2005
R2194 VSS.n1985 VSS.n1984 5.2005
R2195 VSS.n1995 VSS.n1985 5.2005
R2196 VSS.n1993 VSS.n1992 5.2005
R2197 VSS.n1994 VSS.n1993 5.2005
R2198 VSS.n1991 VSS.n1987 5.2005
R2199 VSS.n1987 VSS.n1986 5.2005
R2200 VSS.n1990 VSS.n1989 5.2005
R2201 VSS.n1989 VSS.n1988 5.2005
R2202 VSS.n631 VSS.n630 5.2005
R2203 VSS.n632 VSS.n631 5.2005
R2204 VSS.n2203 VSS.n2202 5.2005
R2205 VSS.n2202 VSS.n2201 5.2005
R2206 VSS.n2206 VSS.n2205 5.2005
R2207 VSS.n2207 VSS.n2206 5.2005
R2208 VSS.n626 VSS.n625 5.2005
R2209 VSS.n2208 VSS.n626 5.2005
R2210 VSS.n2211 VSS.n2210 5.2005
R2211 VSS.n2210 VSS.n2209 5.2005
R2212 VSS.n2212 VSS.n624 5.2005
R2213 VSS.n624 VSS.n623 5.2005
R2214 VSS.n2214 VSS.n2213 5.2005
R2215 VSS.n2215 VSS.n2214 5.2005
R2216 VSS.n622 VSS.n621 5.2005
R2217 VSS.n2216 VSS.n622 5.2005
R2218 VSS.n2219 VSS.n2218 5.2005
R2219 VSS.n2218 VSS.n2217 5.2005
R2220 VSS.n2220 VSS.n620 5.2005
R2221 VSS.n620 VSS.n619 5.2005
R2222 VSS.n2224 VSS.n2223 5.2005
R2223 VSS.n2225 VSS.n2224 5.2005
R2224 VSS.n618 VSS.n617 5.2005
R2225 VSS.n2226 VSS.n618 5.2005
R2226 VSS.n2229 VSS.n2228 5.2005
R2227 VSS.n2228 VSS.n2227 5.2005
R2228 VSS.n2230 VSS.n616 5.2005
R2229 VSS.n616 VSS.n615 5.2005
R2230 VSS.n2232 VSS.n2231 5.2005
R2231 VSS.n2233 VSS.n2232 5.2005
R2232 VSS.n614 VSS.n613 5.2005
R2233 VSS.n2234 VSS.n614 5.2005
R2234 VSS.n2237 VSS.n2236 5.2005
R2235 VSS.n2236 VSS.n2235 5.2005
R2236 VSS.n2238 VSS.n612 5.2005
R2237 VSS.n612 VSS.n611 5.2005
R2238 VSS.n2240 VSS.n2239 5.2005
R2239 VSS.n2241 VSS.n2240 5.2005
R2240 VSS.n610 VSS.n609 5.2005
R2241 VSS.n2242 VSS.n610 5.2005
R2242 VSS.n2245 VSS.n2244 5.2005
R2243 VSS.n2244 VSS.n2243 5.2005
R2244 VSS.n2299 VSS.n2298 5.2005
R2245 VSS.n2298 VSS.n2297 5.2005
R2246 VSS.n2247 VSS.n2246 5.2005
R2247 VSS.n2296 VSS.n2247 5.2005
R2248 VSS.n2294 VSS.n2293 5.2005
R2249 VSS.n2295 VSS.n2294 5.2005
R2250 VSS.n2292 VSS.n2250 5.2005
R2251 VSS.n2250 VSS.n2249 5.2005
R2252 VSS.n2291 VSS.n2290 5.2005
R2253 VSS.n2290 VSS.n2289 5.2005
R2254 VSS.n2252 VSS.n2251 5.2005
R2255 VSS.n2288 VSS.n2252 5.2005
R2256 VSS.n2286 VSS.n2285 5.2005
R2257 VSS.n2287 VSS.n2286 5.2005
R2258 VSS.n2284 VSS.n2254 5.2005
R2259 VSS.n2254 VSS.n2253 5.2005
R2260 VSS.n2283 VSS.n2282 5.2005
R2261 VSS.n2282 VSS.n2281 5.2005
R2262 VSS.n2260 VSS.n2257 5.2005
R2263 VSS.n2280 VSS.n2257 5.2005
R2264 VSS.n2278 VSS.n2277 5.2005
R2265 VSS.n2279 VSS.n2278 5.2005
R2266 VSS.n2276 VSS.n2259 5.2005
R2267 VSS.n2259 VSS.n2258 5.2005
R2268 VSS.n2275 VSS.n2274 5.2005
R2269 VSS.n2274 VSS.n2273 5.2005
R2270 VSS.n2262 VSS.n2261 5.2005
R2271 VSS.n2272 VSS.n2262 5.2005
R2272 VSS.n2270 VSS.n2269 5.2005
R2273 VSS.n2271 VSS.n2270 5.2005
R2274 VSS.n2268 VSS.n2264 5.2005
R2275 VSS.n2264 VSS.n2263 5.2005
R2276 VSS.n2267 VSS.n2266 5.2005
R2277 VSS.n2266 VSS.n2265 5.2005
R2278 VSS.n451 VSS.n450 5.2005
R2279 VSS.n453 VSS.n451 5.2005
R2280 VSS.n2530 VSS.n2529 5.2005
R2281 VSS.n2529 VSS.n2528 5.2005
R2282 VSS.n2532 VSS.n448 5.2005
R2283 VSS.n448 VSS.n447 5.2005
R2284 VSS.n2534 VSS.n2533 5.2005
R2285 VSS.n2535 VSS.n2534 5.2005
R2286 VSS.n446 VSS.n445 5.2005
R2287 VSS.n2536 VSS.n446 5.2005
R2288 VSS.n2539 VSS.n2538 5.2005
R2289 VSS.n2538 VSS.n2537 5.2005
R2290 VSS.n2540 VSS.n444 5.2005
R2291 VSS.n444 VSS.n443 5.2005
R2292 VSS.n2542 VSS.n2541 5.2005
R2293 VSS.n2543 VSS.n2542 5.2005
R2294 VSS.n442 VSS.n441 5.2005
R2295 VSS.n2544 VSS.n442 5.2005
R2296 VSS.n2547 VSS.n2546 5.2005
R2297 VSS.n2546 VSS.n2545 5.2005
R2298 VSS.n2548 VSS.n439 5.2005
R2299 VSS.n439 VSS.n438 5.2005
R2300 VSS.n2551 VSS.n2550 5.2005
R2301 VSS.n2552 VSS.n2551 5.2005
R2302 VSS.n437 VSS.n436 5.2005
R2303 VSS.n2553 VSS.n437 5.2005
R2304 VSS.n2556 VSS.n2555 5.2005
R2305 VSS.n2555 VSS.n2554 5.2005
R2306 VSS.n2557 VSS.n435 5.2005
R2307 VSS.n435 VSS.n434 5.2005
R2308 VSS.n2559 VSS.n2558 5.2005
R2309 VSS.n2560 VSS.n2559 5.2005
R2310 VSS.n433 VSS.n432 5.2005
R2311 VSS.n2561 VSS.n433 5.2005
R2312 VSS.n2565 VSS.n2564 5.2005
R2313 VSS.n2564 VSS.n2563 5.2005
R2314 VSS.n2566 VSS.n431 5.2005
R2315 VSS.n2562 VSS.n431 5.2005
R2316 VSS.n2568 VSS.n2567 5.2005
R2317 VSS.n2568 VSS.n430 5.2005
R2318 VSS.n2569 VSS.n424 5.2005
R2319 VSS.n2570 VSS.n2569 5.2005
R2320 VSS.n2584 VSS.n2583 5.2005
R2321 VSS.n2585 VSS.n2584 5.2005
R2322 VSS.n421 VSS.n420 5.2005
R2323 VSS.n2586 VSS.n421 5.2005
R2324 VSS.n2590 VSS.n2589 5.2005
R2325 VSS.n2589 VSS.n2588 5.2005
R2326 VSS.n2591 VSS.n419 5.2005
R2327 VSS.n2587 VSS.n419 5.2005
R2328 VSS.n2593 VSS.n2592 5.2005
R2329 VSS.n2594 VSS.n2593 5.2005
R2330 VSS.n416 VSS.n415 5.2005
R2331 VSS.n2596 VSS.n416 5.2005
R2332 VSS.n2599 VSS.n2598 5.2005
R2333 VSS.n2598 VSS.n2597 5.2005
R2334 VSS.n2600 VSS.n414 5.2005
R2335 VSS.n414 VSS.n413 5.2005
R2336 VSS.n2603 VSS.n2602 5.2005
R2337 VSS.n2604 VSS.n2603 5.2005
R2338 VSS.n2601 VSS.n412 5.2005
R2339 VSS.n2605 VSS.n412 5.2005
R2340 VSS.n2608 VSS.n2607 5.2005
R2341 VSS.n2607 VSS.n2606 5.2005
R2342 VSS.n2609 VSS.n409 5.2005
R2343 VSS.n409 VSS.n408 5.2005
R2344 VSS.n2611 VSS.n2610 5.2005
R2345 VSS.n2612 VSS.n2611 5.2005
R2346 VSS.n407 VSS.n406 5.2005
R2347 VSS.n2613 VSS.n407 5.2005
R2348 VSS.n2616 VSS.n2615 5.2005
R2349 VSS.n2615 VSS.n2614 5.2005
R2350 VSS.n2617 VSS.n405 5.2005
R2351 VSS.n405 VSS.n404 5.2005
R2352 VSS.n2619 VSS.n2618 5.2005
R2353 VSS.n2620 VSS.n2619 5.2005
R2354 VSS.n402 VSS.n401 5.2005
R2355 VSS.n2621 VSS.n402 5.2005
R2356 VSS.n2654 VSS.n2653 5.2005
R2357 VSS.n2653 VSS.n2652 5.2005
R2358 VSS.n2656 VSS.n399 5.2005
R2359 VSS.n399 VSS.n398 5.2005
R2360 VSS.n2659 VSS.n2658 5.2005
R2361 VSS.n2660 VSS.n2659 5.2005
R2362 VSS.n2657 VSS.n397 5.2005
R2363 VSS.n2661 VSS.n397 5.2005
R2364 VSS.n2663 VSS.n396 5.2005
R2365 VSS.n2663 VSS.n2662 5.2005
R2366 VSS.n2665 VSS.n2664 5.2005
R2367 VSS.n2664 VSS.n392 5.2005
R2368 VSS.n2666 VSS.n393 5.2005
R2369 VSS.n2696 VSS.n2695 5.2005
R2370 VSS.n2697 VSS.n2696 5.2005
R2371 VSS.n2694 VSS.n395 5.2005
R2372 VSS.n395 VSS.n394 5.2005
R2373 VSS.n2693 VSS.n2692 5.2005
R2374 VSS.n2692 VSS.n2691 5.2005
R2375 VSS.n2668 VSS.n2667 5.2005
R2376 VSS.n2690 VSS.n2668 5.2005
R2377 VSS.n2688 VSS.n2687 5.2005
R2378 VSS.n2689 VSS.n2688 5.2005
R2379 VSS.n2686 VSS.n2670 5.2005
R2380 VSS.n2670 VSS.n2669 5.2005
R2381 VSS.n2685 VSS.n2684 5.2005
R2382 VSS.n2684 VSS.n2683 5.2005
R2383 VSS.n2672 VSS.n2671 5.2005
R2384 VSS.n2682 VSS.n2672 5.2005
R2385 VSS.n2680 VSS.n2679 5.2005
R2386 VSS.n2681 VSS.n2680 5.2005
R2387 VSS.n2678 VSS.n2674 5.2005
R2388 VSS.n2674 VSS.n2673 5.2005
R2389 VSS.n2677 VSS.n2676 5.2005
R2390 VSS.n2676 VSS.n2675 5.2005
R2391 VSS.n122 VSS.n121 5.2005
R2392 VSS.n124 VSS.n122 5.2005
R2393 VSS.n3241 VSS.n3240 5.2005
R2394 VSS.n3240 VSS.n3239 5.2005
R2395 VSS.n764 VSS.n715 5.2005
R2396 VSS.n763 VSS.n762 5.2005
R2397 VSS.n761 VSS.n760 5.2005
R2398 VSS.n759 VSS.n758 5.2005
R2399 VSS.n757 VSS.n726 5.2005
R2400 VSS.n741 VSS.n727 5.2005
R2401 VSS.n743 VSS.n742 5.2005
R2402 VSS.n745 VSS.n744 5.2005
R2403 VSS.n747 VSS.n746 5.2005
R2404 VSS.n749 VSS.n748 5.2005
R2405 VSS.n751 VSS.n750 5.2005
R2406 VSS.n752 VSS.n732 5.2005
R2407 VSS.n754 VSS.n753 5.2005
R2408 VSS.n755 VSS.n754 5.2005
R2409 VSS.n349 VSS.n302 5.2005
R2410 VSS.n347 VSS.n346 5.2005
R2411 VSS.n345 VSS.n304 5.2005
R2412 VSS.n344 VSS.n343 5.2005
R2413 VSS.n341 VSS.n305 5.2005
R2414 VSS.n339 VSS.n338 5.2005
R2415 VSS.n337 VSS.n306 5.2005
R2416 VSS.n336 VSS.n335 5.2005
R2417 VSS.n333 VSS.n307 5.2005
R2418 VSS.n333 VSS.n332 5.2005
R2419 VSS.n325 VSS.n308 5.2005
R2420 VSS.n330 VSS.n308 5.2005
R2421 VSS.n327 VSS.n326 5.2005
R2422 VSS.n324 VSS.n309 5.2005
R2423 VSS.n323 VSS.n322 5.2005
R2424 VSS.n322 VSS.n321 5.2005
R2425 VSS.n311 VSS.n310 5.2005
R2426 VSS.n320 VSS.n311 5.2005
R2427 VSS.n318 VSS.n317 5.2005
R2428 VSS.n319 VSS.n318 5.2005
R2429 VSS.n316 VSS.n315 5.2005
R2430 VSS.n315 VSS.n312 5.2005
R2431 VSS.n314 VSS.n153 5.2005
R2432 VSS.n314 VSS.n313 5.2005
R2433 VSS.n2648 VSS.n400 5.2005
R2434 VSS.n2647 VSS.n2646 5.2005
R2435 VSS.n2645 VSS.n2626 5.2005
R2436 VSS.n2644 VSS.n2643 5.2005
R2437 VSS.n2642 VSS.n2641 5.2005
R2438 VSS.n2640 VSS.n2639 5.2005
R2439 VSS.n2638 VSS.n2637 5.2005
R2440 VSS.n2636 VSS.n2632 5.2005
R2441 VSS.n2631 VSS.n2627 5.2005
R2442 VSS.n2631 VSS.n2622 5.2005
R2443 VSS.n2630 VSS.n2628 5.2005
R2444 VSS.n2630 VSS.n2629 5.2005
R2445 VSS.n292 VSS.n291 5.2005
R2446 VSS.n293 VSS.n292 5.2005
R2447 VSS.n2703 VSS.n2702 5.2005
R2448 VSS.n2702 VSS.n2701 5.2005
R2449 VSS.n2704 VSS.n289 5.2005
R2450 VSS.n289 VSS.n287 5.2005
R2451 VSS.n2706 VSS.n2705 5.2005
R2452 VSS.n2707 VSS.n2706 5.2005
R2453 VSS.n290 VSS.n288 5.2005
R2454 VSS.n356 VSS.n353 5.2005
R2455 VSS.n358 VSS.n357 5.2005
R2456 VSS.n359 VSS.n352 5.2005
R2457 VSS.n361 VSS.n360 5.2005
R2458 VSS.n363 VSS.n351 5.2005
R2459 VSS.n364 VSS.n303 5.2005
R2460 VSS.n367 VSS.n366 5.2005
R2461 VSS.n3208 VSS.n3207 5.2005
R2462 VSS.n3209 VSS.n138 5.2005
R2463 VSS.n3211 VSS.n3210 5.2005
R2464 VSS.n3213 VSS.n137 5.2005
R2465 VSS.n3214 VSS.n136 5.2005
R2466 VSS.n3217 VSS.n3216 5.2005
R2467 VSS.n3218 VSS.n134 5.2005
R2468 VSS.n134 VSS.n130 5.2005
R2469 VSS.n3220 VSS.n3219 5.2005
R2470 VSS.n3221 VSS.n3220 5.2005
R2471 VSS.n135 VSS.n133 5.2005
R2472 VSS.n133 VSS.n132 5.2005
R2473 VSS.n381 VSS.n380 5.2005
R2474 VSS.n382 VSS.n381 5.2005
R2475 VSS.n379 VSS.n378 5.2005
R2476 VSS.n383 VSS.n379 5.2005
R2477 VSS.n386 VSS.n385 5.2005
R2478 VSS.n385 VSS.n384 5.2005
R2479 VSS.n387 VSS.n297 5.2005
R2480 VSS.n297 VSS.n295 5.2005
R2481 VSS.n389 VSS.n388 5.2005
R2482 VSS.n390 VSS.n389 5.2005
R2483 VSS.n377 VSS.n296 5.2005
R2484 VSS.n296 VSS.n294 5.2005
R2485 VSS.n376 VSS.n375 5.2005
R2486 VSS.n375 VSS.n374 5.2005
R2487 VSS.n299 VSS.n298 5.2005
R2488 VSS.n373 VSS.n299 5.2005
R2489 VSS.n371 VSS.n370 5.2005
R2490 VSS.n372 VSS.n371 5.2005
R2491 VSS.n369 VSS.n301 5.2005
R2492 VSS.n301 VSS.n300 5.2005
R2493 VSS.n285 VSS.n284 5.2005
R2494 VSS.n2709 VSS.n285 5.2005
R2495 VSS.n2712 VSS.n2711 5.2005
R2496 VSS.n2711 VSS.n2710 5.2005
R2497 VSS.n2713 VSS.n283 5.2005
R2498 VSS.n283 VSS.n282 5.2005
R2499 VSS.n2715 VSS.n2714 5.2005
R2500 VSS.n2716 VSS.n2715 5.2005
R2501 VSS.n281 VSS.n280 5.2005
R2502 VSS.n2717 VSS.n281 5.2005
R2503 VSS.n2720 VSS.n2719 5.2005
R2504 VSS.n2719 VSS.n2718 5.2005
R2505 VSS.n2721 VSS.n279 5.2005
R2506 VSS.n279 VSS.n278 5.2005
R2507 VSS.n2723 VSS.n2722 5.2005
R2508 VSS.n2724 VSS.n2723 5.2005
R2509 VSS.n272 VSS.n271 5.2005
R2510 VSS.n2725 VSS.n272 5.2005
R2511 VSS.n2728 VSS.n2727 5.2005
R2512 VSS.n2727 VSS.n2726 5.2005
R2513 VSS.n2729 VSS.n270 5.2005
R2514 VSS.n276 VSS.n270 5.2005
R2515 VSS.n2731 VSS.n2730 5.2005
R2516 VSS.n2733 VSS.n269 5.2005
R2517 VSS.n2734 VSS.n267 5.2005
R2518 VSS.n2737 VSS.n2736 5.2005
R2519 VSS.n2738 VSS.n266 5.2005
R2520 VSS.n266 VSS.n265 5.2005
R2521 VSS.n2740 VSS.n2739 5.2005
R2522 VSS.n2741 VSS.n2740 5.2005
R2523 VSS.n264 VSS.n263 5.2005
R2524 VSS.n2742 VSS.n264 5.2005
R2525 VSS.n2745 VSS.n2744 5.2005
R2526 VSS.n2744 VSS.n2743 5.2005
R2527 VSS.n2398 VSS.n262 5.2005
R2528 VSS.n2447 VSS.n2398 5.2005
R2529 VSS.n2451 VSS.n2450 5.2005
R2530 VSS.n2450 VSS.n2449 5.2005
R2531 VSS.n2452 VSS.n2397 5.2005
R2532 VSS.n2397 VSS.n2396 5.2005
R2533 VSS.n2454 VSS.n2453 5.2005
R2534 VSS.n2455 VSS.n2454 5.2005
R2535 VSS.n2395 VSS.n2394 5.2005
R2536 VSS.n2456 VSS.n2395 5.2005
R2537 VSS.n2459 VSS.n2458 5.2005
R2538 VSS.n2458 VSS.n2457 5.2005
R2539 VSS.n2460 VSS.n2393 5.2005
R2540 VSS.n2393 VSS.n2392 5.2005
R2541 VSS.n2462 VSS.n2461 5.2005
R2542 VSS.n2463 VSS.n2462 5.2005
R2543 VSS.n2391 VSS.n2390 5.2005
R2544 VSS.n2464 VSS.n2391 5.2005
R2545 VSS.n2467 VSS.n2466 5.2005
R2546 VSS.n2466 VSS.n2465 5.2005
R2547 VSS.n2468 VSS.n2389 5.2005
R2548 VSS.n2389 VSS.n2388 5.2005
R2549 VSS.n2470 VSS.n2469 5.2005
R2550 VSS.n2471 VSS.n2470 5.2005
R2551 VSS.n2387 VSS.n2386 5.2005
R2552 VSS.n2472 VSS.n2387 5.2005
R2553 VSS.n2475 VSS.n2474 5.2005
R2554 VSS.n2474 VSS.n2473 5.2005
R2555 VSS.n2476 VSS.n2384 5.2005
R2556 VSS.n2384 VSS.n2383 5.2005
R2557 VSS.n2478 VSS.n2477 5.2005
R2558 VSS.n2479 VSS.n2478 5.2005
R2559 VSS.n2385 VSS.n2382 5.2005
R2560 VSS.n2480 VSS.n2382 5.2005
R2561 VSS.n2482 VSS.n2381 5.2005
R2562 VSS.n2482 VSS.n2481 5.2005
R2563 VSS.n2484 VSS.n2483 5.2005
R2564 VSS.n2483 VSS.n192 5.2005
R2565 VSS.n2380 VSS.n2379 5.2005
R2566 VSS.n2379 VSS.n474 5.2005
R2567 VSS.n2378 VSS.n518 5.2005
R2568 VSS.n2378 VSS.n2377 5.2005
R2569 VSS.n2372 VSS.n519 5.2005
R2570 VSS.n2376 VSS.n519 5.2005
R2571 VSS.n2374 VSS.n2373 5.2005
R2572 VSS.n2375 VSS.n2374 5.2005
R2573 VSS.n2371 VSS.n521 5.2005
R2574 VSS.n521 VSS.n520 5.2005
R2575 VSS.n2370 VSS.n2369 5.2005
R2576 VSS.n2369 VSS.n2368 5.2005
R2577 VSS.n523 VSS.n522 5.2005
R2578 VSS.n2367 VSS.n523 5.2005
R2579 VSS.n2365 VSS.n2364 5.2005
R2580 VSS.n2366 VSS.n2365 5.2005
R2581 VSS.n2363 VSS.n525 5.2005
R2582 VSS.n525 VSS.n524 5.2005
R2583 VSS.n2362 VSS.n2361 5.2005
R2584 VSS.n2361 VSS.n2360 5.2005
R2585 VSS.n527 VSS.n526 5.2005
R2586 VSS.n2359 VSS.n527 5.2005
R2587 VSS.n2357 VSS.n2356 5.2005
R2588 VSS.n2358 VSS.n2357 5.2005
R2589 VSS.n2355 VSS.n529 5.2005
R2590 VSS.n529 VSS.n528 5.2005
R2591 VSS.n2354 VSS.n2353 5.2005
R2592 VSS.n2353 VSS.n2352 5.2005
R2593 VSS.n531 VSS.n530 5.2005
R2594 VSS.n2351 VSS.n531 5.2005
R2595 VSS.n2349 VSS.n2348 5.2005
R2596 VSS.n2350 VSS.n2349 5.2005
R2597 VSS.n2347 VSS.n533 5.2005
R2598 VSS.n533 VSS.n532 5.2005
R2599 VSS.n2346 VSS.n2345 5.2005
R2600 VSS.n2345 VSS.n2344 5.2005
R2601 VSS.n2342 VSS.n534 5.2005
R2602 VSS.n2343 VSS.n2342 5.2005
R2603 VSS.n2340 VSS.n538 5.2005
R2604 VSS.n2340 VSS.n2339 5.2005
R2605 VSS.n2119 VSS.n537 5.2005
R2606 VSS.n539 VSS.n537 5.2005
R2607 VSS.n2122 VSS.n2121 5.2005
R2608 VSS.n2121 VSS.n2120 5.2005
R2609 VSS.n2123 VSS.n2118 5.2005
R2610 VSS.n2118 VSS.n2117 5.2005
R2611 VSS.n2125 VSS.n2124 5.2005
R2612 VSS.n2126 VSS.n2125 5.2005
R2613 VSS.n2116 VSS.n2115 5.2005
R2614 VSS.n2127 VSS.n2116 5.2005
R2615 VSS.n2130 VSS.n2129 5.2005
R2616 VSS.n2129 VSS.n2128 5.2005
R2617 VSS.n2131 VSS.n2114 5.2005
R2618 VSS.n2114 VSS.n2113 5.2005
R2619 VSS.n2133 VSS.n2132 5.2005
R2620 VSS.n2134 VSS.n2133 5.2005
R2621 VSS.n2112 VSS.n2111 5.2005
R2622 VSS.n2135 VSS.n2112 5.2005
R2623 VSS.n2138 VSS.n2137 5.2005
R2624 VSS.n2137 VSS.n2136 5.2005
R2625 VSS.n2139 VSS.n2110 5.2005
R2626 VSS.n2110 VSS.n2109 5.2005
R2627 VSS.n2141 VSS.n2140 5.2005
R2628 VSS.n2142 VSS.n2141 5.2005
R2629 VSS.n2108 VSS.n2107 5.2005
R2630 VSS.n2143 VSS.n2108 5.2005
R2631 VSS.n2146 VSS.n2145 5.2005
R2632 VSS.n2145 VSS.n2144 5.2005
R2633 VSS.n2147 VSS.n2106 5.2005
R2634 VSS.n2106 VSS.n2105 5.2005
R2635 VSS.n2149 VSS.n2148 5.2005
R2636 VSS.n2150 VSS.n2149 5.2005
R2637 VSS.n2104 VSS.n695 5.2005
R2638 VSS.n2151 VSS.n2104 5.2005
R2639 VSS.n2154 VSS.n2153 5.2005
R2640 VSS.n2153 VSS.n2152 5.2005
R2641 VSS.n2102 VSS.n694 5.2005
R2642 VSS.n2102 VSS.n649 5.2005
R2643 VSS.n2101 VSS.n698 5.2005
R2644 VSS.n2101 VSS.n2100 5.2005
R2645 VSS.n2095 VSS.n697 5.2005
R2646 VSS.n2099 VSS.n697 5.2005
R2647 VSS.n2097 VSS.n2096 5.2005
R2648 VSS.n2098 VSS.n2097 5.2005
R2649 VSS.n2094 VSS.n700 5.2005
R2650 VSS.n700 VSS.n699 5.2005
R2651 VSS.n2093 VSS.n2092 5.2005
R2652 VSS.n2092 VSS.n2091 5.2005
R2653 VSS.n702 VSS.n701 5.2005
R2654 VSS.n2090 VSS.n702 5.2005
R2655 VSS.n2088 VSS.n2087 5.2005
R2656 VSS.n2089 VSS.n2088 5.2005
R2657 VSS.n2086 VSS.n704 5.2005
R2658 VSS.n704 VSS.n703 5.2005
R2659 VSS.n2085 VSS.n2084 5.2005
R2660 VSS.n2084 VSS.n2083 5.2005
R2661 VSS.n706 VSS.n705 5.2005
R2662 VSS.n2082 VSS.n706 5.2005
R2663 VSS.n2080 VSS.n2079 5.2005
R2664 VSS.n2081 VSS.n2080 5.2005
R2665 VSS.n2078 VSS.n708 5.2005
R2666 VSS.n708 VSS.n707 5.2005
R2667 VSS.n2077 VSS.n2076 5.2005
R2668 VSS.n2076 VSS.n2075 5.2005
R2669 VSS.n710 VSS.n709 5.2005
R2670 VSS.n2074 VSS.n710 5.2005
R2671 VSS.n2072 VSS.n2071 5.2005
R2672 VSS.n2073 VSS.n2072 5.2005
R2673 VSS.n2070 VSS.n712 5.2005
R2674 VSS.n712 VSS.n711 5.2005
R2675 VSS.n2069 VSS.n2068 5.2005
R2676 VSS.n2068 VSS.n2067 5.2005
R2677 VSS.n2065 VSS.n713 5.2005
R2678 VSS.n2066 VSS.n2065 5.2005
R2679 VSS.n2063 VSS.n717 5.2005
R2680 VSS.n2063 VSS.n2062 5.2005
R2681 VSS.n852 VSS.n716 5.2005
R2682 VSS.n718 VSS.n716 5.2005
R2683 VSS.n855 VSS.n854 5.2005
R2684 VSS.n854 VSS.n853 5.2005
R2685 VSS.n856 VSS.n851 5.2005
R2686 VSS.n851 VSS.n850 5.2005
R2687 VSS.n858 VSS.n857 5.2005
R2688 VSS.n859 VSS.n858 5.2005
R2689 VSS.n849 VSS.n848 5.2005
R2690 VSS.n860 VSS.n849 5.2005
R2691 VSS.n863 VSS.n862 5.2005
R2692 VSS.n862 VSS.n861 5.2005
R2693 VSS.n864 VSS.n847 5.2005
R2694 VSS.n847 VSS.n846 5.2005
R2695 VSS.n866 VSS.n865 5.2005
R2696 VSS.n867 VSS.n866 5.2005
R2697 VSS.n845 VSS.n844 5.2005
R2698 VSS.n868 VSS.n845 5.2005
R2699 VSS.n871 VSS.n870 5.2005
R2700 VSS.n870 VSS.n869 5.2005
R2701 VSS.n872 VSS.n843 5.2005
R2702 VSS.n843 VSS.n842 5.2005
R2703 VSS.n874 VSS.n873 5.2005
R2704 VSS.n875 VSS.n874 5.2005
R2705 VSS.n841 VSS.n840 5.2005
R2706 VSS.n876 VSS.n841 5.2005
R2707 VSS.n879 VSS.n878 5.2005
R2708 VSS.n878 VSS.n877 5.2005
R2709 VSS.n880 VSS.n838 5.2005
R2710 VSS.n838 VSS.n837 5.2005
R2711 VSS.n882 VSS.n881 5.2005
R2712 VSS.n883 VSS.n882 5.2005
R2713 VSS.n839 VSS.n835 5.2005
R2714 VSS.n884 VSS.n835 5.2005
R2715 VSS.n886 VSS.n836 5.2005
R2716 VSS.n886 VSS.n885 5.2005
R2717 VSS.n1748 VSS.n834 5.2005
R2718 VSS.n834 VSS.n828 5.2005
R2719 VSS.n1750 VSS.n1749 5.2005
R2720 VSS.n1751 VSS.n1750 5.2005
R2721 VSS.n1747 VSS.n1746 5.2005
R2722 VSS.n1752 VSS.n1747 5.2005
R2723 VSS.n1755 VSS.n1754 5.2005
R2724 VSS.n1754 VSS.n1753 5.2005
R2725 VSS.n1756 VSS.n1745 5.2005
R2726 VSS.n1745 VSS.n1744 5.2005
R2727 VSS.n1758 VSS.n1757 5.2005
R2728 VSS.n1759 VSS.n1758 5.2005
R2729 VSS.n1743 VSS.n1742 5.2005
R2730 VSS.n1760 VSS.n1743 5.2005
R2731 VSS.n1763 VSS.n1762 5.2005
R2732 VSS.n1762 VSS.n1761 5.2005
R2733 VSS.n1764 VSS.n1741 5.2005
R2734 VSS.n1741 VSS.n1740 5.2005
R2735 VSS.n1766 VSS.n1765 5.2005
R2736 VSS.n1767 VSS.n1766 5.2005
R2737 VSS.n1739 VSS.n1738 5.2005
R2738 VSS.n1768 VSS.n1739 5.2005
R2739 VSS.n1771 VSS.n1770 5.2005
R2740 VSS.n1770 VSS.n1769 5.2005
R2741 VSS.n1772 VSS.n1736 5.2005
R2742 VSS.n1736 VSS.n1735 5.2005
R2743 VSS.n1774 VSS.n1773 5.2005
R2744 VSS.n1775 VSS.n1774 5.2005
R2745 VSS.n1737 VSS.n1734 5.2005
R2746 VSS.n1776 VSS.n1734 5.2005
R2747 VSS.n1778 VSS.n1733 5.2005
R2748 VSS.n1778 VSS.n1777 5.2005
R2749 VSS.n1780 VSS.n1779 5.2005
R2750 VSS.n1779 VSS.n890 5.2005
R2751 VSS.n1781 VSS.n918 5.2005
R2752 VSS.n918 VSS.n916 5.2005
R2753 VSS.n1783 VSS.n1782 5.2005
R2754 VSS.n1784 VSS.n1783 5.2005
R2755 VSS.n1876 VSS.n1875 5.2005
R2756 VSS.n1874 VSS.n1873 5.2005
R2757 VSS.n1872 VSS.n1871 5.2005
R2758 VSS.n1870 VSS.n1869 5.2005
R2759 VSS.n1868 VSS.n887 5.2005
R2760 VSS.n1852 VSS.n888 5.2005
R2761 VSS.n1854 VSS.n1853 5.2005
R2762 VSS.n1856 VSS.n1855 5.2005
R2763 VSS.n1858 VSS.n1857 5.2005
R2764 VSS.n1860 VSS.n1859 5.2005
R2765 VSS.n1862 VSS.n1861 5.2005
R2766 VSS.n1863 VSS.n1842 5.2005
R2767 VSS.n1865 VSS.n1864 5.2005
R2768 VSS.n1866 VSS.n1865 5.2005
R2769 VSS.n1788 VSS.n1787 5.2005
R2770 VSS.n911 VSS.n910 5.2005
R2771 VSS.n921 VSS.n920 5.2005
R2772 VSS.n923 VSS.n922 5.2005
R2773 VSS.n1730 VSS.n1729 5.2005
R2774 VSS.n1728 VSS.n1727 5.2005
R2775 VSS.n925 VSS.n924 5.2005
R2776 VSS.n1589 VSS.n1588 5.2005
R2777 VSS.n1592 VSS.n1591 5.2005
R2778 VSS.n1591 VSS.n1590 5.2005
R2779 VSS.n1593 VSS.n1587 5.2005
R2780 VSS.n1587 VSS.n1586 5.2005
R2781 VSS.n1595 VSS.n1594 5.2005
R2782 VSS.n1596 VSS.n1595 5.2005
R2783 VSS.n1585 VSS.n1584 5.2005
R2784 VSS.n1597 VSS.n1585 5.2005
R2785 VSS.n1601 VSS.n1600 5.2005
R2786 VSS.n1600 VSS.n1599 5.2005
R2787 VSS.n1602 VSS.n1583 5.2005
R2788 VSS.n1598 VSS.n1583 5.2005
R2789 VSS.n1604 VSS.n1603 5.2005
R2790 VSS.n1604 VSS.n1567 5.2005
R2791 VSS.n1606 VSS.n1605 5.2005
R2792 VSS.n1605 VSS.n1568 5.2005
R2793 VSS.n1607 VSS.n1582 5.2005
R2794 VSS.n1582 VSS.n1581 5.2005
R2795 VSS.n1609 VSS.n1608 5.2005
R2796 VSS.n1610 VSS.n1609 5.2005
R2797 VSS.n1580 VSS.n1579 5.2005
R2798 VSS.n1611 VSS.n1580 5.2005
R2799 VSS.n1614 VSS.n1613 5.2005
R2800 VSS.n1613 VSS.n1612 5.2005
R2801 VSS.n1615 VSS.n1577 5.2005
R2802 VSS.n1577 VSS.n1576 5.2005
R2803 VSS.n1624 VSS.n1623 5.2005
R2804 VSS.n1625 VSS.n1624 5.2005
R2805 VSS.n1622 VSS.n1578 5.2005
R2806 VSS.n1621 VSS.n1620 5.2005
R2807 VSS.n1619 VSS.n1618 5.2005
R2808 VSS.n1617 VSS.n1616 5.2005
R2809 VSS.n1490 VSS.n1489 5.2005
R2810 VSS.n1489 VSS.n1488 5.2005
R2811 VSS.n1065 VSS.n1064 5.2005
R2812 VSS.n1487 VSS.n1065 5.2005
R2813 VSS.n1485 VSS.n1484 5.2005
R2814 VSS.n1486 VSS.n1485 5.2005
R2815 VSS.n1483 VSS.n1067 5.2005
R2816 VSS.n1067 VSS.n1066 5.2005
R2817 VSS.n1482 VSS.n1481 5.2005
R2818 VSS.n1481 VSS.n1480 5.2005
R2819 VSS.n1069 VSS.n1068 5.2005
R2820 VSS.n1479 VSS.n1069 5.2005
R2821 VSS.n1477 VSS.n1476 5.2005
R2822 VSS.n1478 VSS.n1477 5.2005
R2823 VSS.n1475 VSS.n1071 5.2005
R2824 VSS.n1071 VSS.n1070 5.2005
R2825 VSS.n1513 VSS.n1512 5.2005
R2826 VSS.n1512 VSS.n1511 5.2005
R2827 VSS.n1008 VSS.n1007 5.2005
R2828 VSS.n1509 VSS.n1008 5.2005
R2829 VSS.n1507 VSS.n1506 5.2005
R2830 VSS.n1508 VSS.n1507 5.2005
R2831 VSS.n1505 VSS.n1010 5.2005
R2832 VSS.n1010 VSS.n1009 5.2005
R2833 VSS.n1504 VSS.n1503 5.2005
R2834 VSS.n1503 VSS.n1502 5.2005
R2835 VSS.n1012 VSS.n1011 5.2005
R2836 VSS.n1501 VSS.n1012 5.2005
R2837 VSS.n1499 VSS.n1498 5.2005
R2838 VSS.n1500 VSS.n1499 5.2005
R2839 VSS.n1181 VSS.n1180 5.2005
R2840 VSS.n1183 VSS.n1182 5.2005
R2841 VSS.n1115 VSS.n1106 5.2005
R2842 VSS.n1117 VSS.n1116 5.2005
R2843 VSS.n1116 VSS.n1104 5.2005
R2844 VSS.n1124 VSS.n1096 5.2005
R2845 VSS.n1125 VSS.n1095 5.2005
R2846 VSS.n1198 VSS.n1095 5.2005
R2847 VSS.n1127 VSS.n1126 5.2005
R2848 VSS.n1129 VSS.n1128 5.2005
R2849 VSS.n1131 VSS.n1130 5.2005
R2850 VSS.n1133 VSS.n1132 5.2005
R2851 VSS.n1135 VSS.n1134 5.2005
R2852 VSS.n1137 VSS.n1136 5.2005
R2853 VSS.n1139 VSS.n1138 5.2005
R2854 VSS.n1141 VSS.n1140 5.2005
R2855 VSS.n1143 VSS.n1142 5.2005
R2856 VSS.n1145 VSS.n1144 5.2005
R2857 VSS.n1147 VSS.n1146 5.2005
R2858 VSS.n1149 VSS.n1148 5.2005
R2859 VSS.n1151 VSS.n1150 5.2005
R2860 VSS.n1155 VSS.n1154 5.2005
R2861 VSS.n1034 VSS.n1033 5.2005
R2862 VSS.n1035 VSS.n1031 5.2005
R2863 VSS.n1037 VSS.n1036 5.2005
R2864 VSS.n1039 VSS.n1029 5.2005
R2865 VSS.n1041 VSS.n1040 5.2005
R2866 VSS.n1042 VSS.n1028 5.2005
R2867 VSS.n1044 VSS.n1043 5.2005
R2868 VSS.n1046 VSS.n1026 5.2005
R2869 VSS.n1048 VSS.n1047 5.2005
R2870 VSS.n1049 VSS.n1025 5.2005
R2871 VSS.n1051 VSS.n1050 5.2005
R2872 VSS.n1053 VSS.n1023 5.2005
R2873 VSS.n1055 VSS.n1054 5.2005
R2874 VSS.n1056 VSS.n1022 5.2005
R2875 VSS.n1058 VSS.n1057 5.2005
R2876 VSS.n1060 VSS.n1021 5.2005
R2877 VSS.n1062 VSS.n1061 5.2005
R2878 VSS.n1061 VSS.n1017 5.2005
R2879 VSS.n1497 VSS.n1014 5.2005
R2880 VSS.n1018 VSS.n1014 5.2005
R2881 VSS.n1496 VSS.n1495 5.2005
R2882 VSS.n1495 VSS.n1494 5.2005
R2883 VSS.n1169 VSS.n1168 5.2005
R2884 VSS.n1170 VSS.n1169 5.2005
R2885 VSS.n1167 VSS.n1122 5.2005
R2886 VSS.n1171 VSS.n1122 5.2005
R2887 VSS.n1166 VSS.n1165 5.2005
R2888 VSS.n1165 VSS.n1121 5.2005
R2889 VSS.n1164 VSS.n1111 5.2005
R2890 VSS.n1177 VSS.n1111 5.2005
R2891 VSS.n1163 VSS.n1110 5.2005
R2892 VSS.n1178 VSS.n1110 5.2005
R2893 VSS.n1162 VSS.n1107 5.2005
R2894 VSS.n1184 VSS.n1107 5.2005
R2895 VSS.n1161 VSS.n1103 5.2005
R2896 VSS.n1188 VSS.n1103 5.2005
R2897 VSS.n1160 VSS.n1102 5.2005
R2898 VSS.n1189 VSS.n1102 5.2005
R2899 VSS.n1159 VSS.n1101 5.2005
R2900 VSS.n1190 VSS.n1101 5.2005
R2901 VSS.n1158 VSS.n1157 5.2005
R2902 VSS.n1157 VSS.n1100 5.2005
R2903 VSS.n1156 VSS.n1123 5.2005
R2904 VSS.n1156 VSS.n1094 5.2005
R2905 VSS.n1195 VSS.n1194 5.2005
R2906 VSS.n1195 VSS.n1094 5.2005
R2907 VSS.n1193 VSS.n1097 5.2005
R2908 VSS.n1100 VSS.n1097 5.2005
R2909 VSS.n1192 VSS.n1191 5.2005
R2910 VSS.n1191 VSS.n1190 5.2005
R2911 VSS.n1099 VSS.n1098 5.2005
R2912 VSS.n1189 VSS.n1099 5.2005
R2913 VSS.n1188 VSS.n1187 5.2005
R2914 VSS.n1185 VSS.n1184 5.2005
R2915 VSS.n1105 VSS.n1072 5.2005
R2916 VSS.n1178 VSS.n1105 5.2005
R2917 VSS.n1176 VSS.n1175 5.2005
R2918 VSS.n1177 VSS.n1176 5.2005
R2919 VSS.n1174 VSS.n1113 5.2005
R2920 VSS.n1121 VSS.n1113 5.2005
R2921 VSS.n1173 VSS.n1172 5.2005
R2922 VSS.n1172 VSS.n1171 5.2005
R2923 VSS.n1120 VSS.n1119 5.2005
R2924 VSS.n1170 VSS.n1120 5.2005
R2925 VSS.n1493 VSS.n1492 5.2005
R2926 VSS.n1494 VSS.n1493 5.2005
R2927 VSS.n1491 VSS.n1020 5.2005
R2928 VSS.n1020 VSS.n1018 5.2005
R2929 VSS.n1514 VSS.n1006 5.2005
R2930 VSS.n1806 VSS.n902 5.2005
R2931 VSS.n1804 VSS.n1803 5.2005
R2932 VSS.n1802 VSS.n903 5.2005
R2933 VSS.n1801 VSS.n1800 5.2005
R2934 VSS.n1798 VSS.n1797 5.2005
R2935 VSS.n1795 VSS.n1794 5.2005
R2936 VSS.n1793 VSS.n908 5.2005
R2937 VSS.n1791 VSS.n1790 5.2005
R2938 VSS.n1789 VSS.n909 5.2005
R2939 VSS.n909 VSS.n891 5.2005
R2940 VSS.n1813 VSS.n1812 5.2005
R2941 VSS.n1811 VSS.n900 5.2005
R2942 VSS.n1810 VSS.n1809 5.2005
R2943 VSS.n1808 VSS.n1807 5.2005
R2944 VSS.n1851 VSS.n1841 5.2005
R2945 VSS.n1850 VSS.n1849 5.2005
R2946 VSS.n1844 VSS.n1843 5.2005
R2947 VSS.n1845 VSS.n19 5.2005
R2948 VSS.n740 VSS.n731 5.2005
R2949 VSS.n739 VSS.n738 5.2005
R2950 VSS.n736 VSS.n733 5.2005
R2951 VSS.n734 VSS.n42 5.2005
R2952 VSS.n669 VSS.n660 5.2005
R2953 VSS.n668 VSS.n667 5.2005
R2954 VSS.n665 VSS.n662 5.2005
R2955 VSS.n663 VSS.n64 5.2005
R2956 VSS.n561 VSS.n552 5.2005
R2957 VSS.n560 VSS.n559 5.2005
R2958 VSS.n557 VSS.n554 5.2005
R2959 VSS.n555 VSS.n86 5.2005
R2960 VSS.n491 VSS.n490 5.2005
R2961 VSS.n489 VSS.n488 5.2005
R2962 VSS.n487 VSS.n486 5.2005
R2963 VSS.n485 VSS.n484 5.2005
R2964 VSS.n2771 VSS.n2770 5.2005
R2965 VSS.n249 VSS.n243 5.2005
R2966 VSS.n248 VSS.n247 5.2005
R2967 VSS.n246 VSS.n245 5.2005
R2968 VSS.n1518 VSS.n1517 5.2005
R2969 VSS.n1520 VSS.n1519 5.2005
R2970 VSS.n1522 VSS.n1521 5.2005
R2971 VSS.n1524 VSS.n1523 5.2005
R2972 VSS.n1526 VSS.n1525 5.2005
R2973 VSS.n1528 VSS.n1527 5.2005
R2974 VSS.n1530 VSS.n1529 5.2005
R2975 VSS.n1532 VSS.n1531 5.2005
R2976 VSS.n1534 VSS.n1533 5.2005
R2977 VSS.n1536 VSS.n1535 5.2005
R2978 VSS.n1538 VSS.n1537 5.2005
R2979 VSS.n1540 VSS.n1539 5.2005
R2980 VSS.n1542 VSS.n1541 5.2005
R2981 VSS.n1544 VSS.n1543 5.2005
R2982 VSS.n1546 VSS.n1545 5.2005
R2983 VSS.n1547 VSS.n1003 5.2005
R2984 VSS.n1549 VSS.n1548 5.2005
R2985 VSS.n1550 VSS.n1549 5.2005
R2986 VSS.n1516 VSS.n1515 5.2005
R2987 VSS.n1516 VSS.n993 5.2005
R2988 VSS.n1474 VSS.n1002 5.2005
R2989 VSS.n1002 VSS.n993 5.2005
R2990 VSS.n1818 VSS.n1817 5.2005
R2991 VSS.n1817 VSS.n1816 5.2005
R2992 VSS.n1819 VSS.n894 5.2005
R2993 VSS.n894 VSS.n892 5.2005
R2994 VSS.n1835 VSS.n1834 5.2005
R2995 VSS.n1836 VSS.n1835 5.2005
R2996 VSS.n1833 VSS.n895 5.2005
R2997 VSS.n895 VSS.n893 5.2005
R2998 VSS.n1832 VSS.n1831 5.2005
R2999 VSS.n1831 VSS.n1830 5.2005
R3000 VSS.n1821 VSS.n1820 5.2005
R3001 VSS.n1829 VSS.n1821 5.2005
R3002 VSS.n1827 VSS.n1826 5.2005
R3003 VSS.n1828 VSS.n1827 5.2005
R3004 VSS.n1825 VSS.n1824 5.2005
R3005 VSS.n1824 VSS.n1822 5.2005
R3006 VSS.n1823 VSS.n7 5.2005
R3007 VSS.n1823 VSS.n4 5.2005
R3008 VSS.n3425 VSS.n3424 5.2005
R3009 VSS.n3425 VSS.n5 5.2005
R3010 VSS.n3422 VSS.n6 5.2005
R3011 VSS.n12 VSS.n6 5.2005
R3012 VSS.n3421 VSS.n3420 5.2005
R3013 VSS.n3420 VSS.n3419 5.2005
R3014 VSS.n11 VSS.n10 5.2005
R3015 VSS.n3418 VSS.n11 5.2005
R3016 VSS.n3416 VSS.n3415 5.2005
R3017 VSS.n3417 VSS.n3416 5.2005
R3018 VSS.n3414 VSS.n14 5.2005
R3019 VSS.n14 VSS.n13 5.2005
R3020 VSS.n3413 VSS.n3412 5.2005
R3021 VSS.n3412 VSS.n3411 5.2005
R3022 VSS.n16 VSS.n15 5.2005
R3023 VSS.n3410 VSS.n16 5.2005
R3024 VSS.n3408 VSS.n3407 5.2005
R3025 VSS.n3409 VSS.n3408 5.2005
R3026 VSS.n3406 VSS.n18 5.2005
R3027 VSS.n18 VSS.n17 5.2005
R3028 VSS.n3404 VSS.n3403 5.2005
R3029 VSS.n3403 VSS.n3402 5.2005
R3030 VSS.n22 VSS.n20 5.2005
R3031 VSS.n3401 VSS.n22 5.2005
R3032 VSS.n3399 VSS.n3398 5.2005
R3033 VSS.n3400 VSS.n3399 5.2005
R3034 VSS.n3397 VSS.n25 5.2005
R3035 VSS.n25 VSS.n24 5.2005
R3036 VSS.n3396 VSS.n3395 5.2005
R3037 VSS.n3395 VSS.n3394 5.2005
R3038 VSS.n27 VSS.n26 5.2005
R3039 VSS.n3393 VSS.n27 5.2005
R3040 VSS.n3391 VSS.n3390 5.2005
R3041 VSS.n3392 VSS.n3391 5.2005
R3042 VSS.n3389 VSS.n29 5.2005
R3043 VSS.n29 VSS.n28 5.2005
R3044 VSS.n3388 VSS.n3387 5.2005
R3045 VSS.n3387 VSS.n3386 5.2005
R3046 VSS.n31 VSS.n30 5.2005
R3047 VSS.n3385 VSS.n31 5.2005
R3048 VSS.n3383 VSS.n3382 5.2005
R3049 VSS.n3384 VSS.n3383 5.2005
R3050 VSS.n3381 VSS.n33 5.2005
R3051 VSS.n33 VSS.n32 5.2005
R3052 VSS.n3380 VSS.n3379 5.2005
R3053 VSS.n3379 VSS.n3378 5.2005
R3054 VSS.n35 VSS.n34 5.2005
R3055 VSS.n3377 VSS.n35 5.2005
R3056 VSS.n3375 VSS.n3374 5.2005
R3057 VSS.n3376 VSS.n3375 5.2005
R3058 VSS.n3373 VSS.n37 5.2005
R3059 VSS.n37 VSS.n36 5.2005
R3060 VSS.n3372 VSS.n3371 5.2005
R3061 VSS.n3371 VSS.n3370 5.2005
R3062 VSS.n39 VSS.n38 5.2005
R3063 VSS.n3369 VSS.n39 5.2005
R3064 VSS.n3367 VSS.n3366 5.2005
R3065 VSS.n3368 VSS.n3367 5.2005
R3066 VSS.n3364 VSS.n3363 5.2005
R3067 VSS.n3363 VSS.n3362 5.2005
R3068 VSS.n44 VSS.n43 5.2005
R3069 VSS.n3361 VSS.n44 5.2005
R3070 VSS.n3359 VSS.n3358 5.2005
R3071 VSS.n3360 VSS.n3359 5.2005
R3072 VSS.n3357 VSS.n47 5.2005
R3073 VSS.n47 VSS.n46 5.2005
R3074 VSS.n3356 VSS.n3355 5.2005
R3075 VSS.n3355 VSS.n3354 5.2005
R3076 VSS.n49 VSS.n48 5.2005
R3077 VSS.n3353 VSS.n49 5.2005
R3078 VSS.n3351 VSS.n3350 5.2005
R3079 VSS.n3352 VSS.n3351 5.2005
R3080 VSS.n3349 VSS.n51 5.2005
R3081 VSS.n51 VSS.n50 5.2005
R3082 VSS.n3348 VSS.n3347 5.2005
R3083 VSS.n3347 VSS.n3346 5.2005
R3084 VSS.n53 VSS.n52 5.2005
R3085 VSS.n3345 VSS.n53 5.2005
R3086 VSS.n3343 VSS.n3342 5.2005
R3087 VSS.n3344 VSS.n3343 5.2005
R3088 VSS.n3341 VSS.n55 5.2005
R3089 VSS.n55 VSS.n54 5.2005
R3090 VSS.n3340 VSS.n3339 5.2005
R3091 VSS.n3339 VSS.n3338 5.2005
R3092 VSS.n57 VSS.n56 5.2005
R3093 VSS.n3337 VSS.n57 5.2005
R3094 VSS.n3335 VSS.n3334 5.2005
R3095 VSS.n3336 VSS.n3335 5.2005
R3096 VSS.n3333 VSS.n59 5.2005
R3097 VSS.n59 VSS.n58 5.2005
R3098 VSS.n3332 VSS.n3331 5.2005
R3099 VSS.n3331 VSS.n3330 5.2005
R3100 VSS.n61 VSS.n60 5.2005
R3101 VSS.n3329 VSS.n61 5.2005
R3102 VSS.n3327 VSS.n3326 5.2005
R3103 VSS.n3328 VSS.n3327 5.2005
R3104 VSS.n3324 VSS.n3323 5.2005
R3105 VSS.n3323 VSS.n3322 5.2005
R3106 VSS.n66 VSS.n65 5.2005
R3107 VSS.n3321 VSS.n66 5.2005
R3108 VSS.n3319 VSS.n3318 5.2005
R3109 VSS.n3320 VSS.n3319 5.2005
R3110 VSS.n3317 VSS.n69 5.2005
R3111 VSS.n69 VSS.n68 5.2005
R3112 VSS.n3316 VSS.n3315 5.2005
R3113 VSS.n3315 VSS.n3314 5.2005
R3114 VSS.n71 VSS.n70 5.2005
R3115 VSS.n3313 VSS.n71 5.2005
R3116 VSS.n3311 VSS.n3310 5.2005
R3117 VSS.n3312 VSS.n3311 5.2005
R3118 VSS.n3309 VSS.n73 5.2005
R3119 VSS.n73 VSS.n72 5.2005
R3120 VSS.n3308 VSS.n3307 5.2005
R3121 VSS.n3307 VSS.n3306 5.2005
R3122 VSS.n75 VSS.n74 5.2005
R3123 VSS.n3305 VSS.n75 5.2005
R3124 VSS.n3303 VSS.n3302 5.2005
R3125 VSS.n3304 VSS.n3303 5.2005
R3126 VSS.n3301 VSS.n77 5.2005
R3127 VSS.n77 VSS.n76 5.2005
R3128 VSS.n3300 VSS.n3299 5.2005
R3129 VSS.n3299 VSS.n3298 5.2005
R3130 VSS.n79 VSS.n78 5.2005
R3131 VSS.n3297 VSS.n79 5.2005
R3132 VSS.n3295 VSS.n3294 5.2005
R3133 VSS.n3296 VSS.n3295 5.2005
R3134 VSS.n3293 VSS.n81 5.2005
R3135 VSS.n81 VSS.n80 5.2005
R3136 VSS.n3292 VSS.n3291 5.2005
R3137 VSS.n3291 VSS.n3290 5.2005
R3138 VSS.n83 VSS.n82 5.2005
R3139 VSS.n3289 VSS.n83 5.2005
R3140 VSS.n3287 VSS.n3286 5.2005
R3141 VSS.n3288 VSS.n3287 5.2005
R3142 VSS.n3284 VSS.n3283 5.2005
R3143 VSS.n3283 VSS.n3282 5.2005
R3144 VSS.n88 VSS.n87 5.2005
R3145 VSS.n3281 VSS.n88 5.2005
R3146 VSS.n3279 VSS.n3278 5.2005
R3147 VSS.n3280 VSS.n3279 5.2005
R3148 VSS.n3277 VSS.n91 5.2005
R3149 VSS.n91 VSS.n90 5.2005
R3150 VSS.n3276 VSS.n3275 5.2005
R3151 VSS.n3275 VSS.n3274 5.2005
R3152 VSS.n93 VSS.n92 5.2005
R3153 VSS.n3273 VSS.n93 5.2005
R3154 VSS.n3271 VSS.n3270 5.2005
R3155 VSS.n3272 VSS.n3271 5.2005
R3156 VSS.n3269 VSS.n94 5.2005
R3157 VSS.n97 VSS.n94 5.2005
R3158 VSS.n3268 VSS.n3267 5.2005
R3159 VSS.n3267 VSS.n3266 5.2005
R3160 VSS.n96 VSS.n95 5.2005
R3161 VSS.n3265 VSS.n96 5.2005
R3162 VSS.n205 VSS.n204 5.2005
R3163 VSS.n204 VSS.n101 5.2005
R3164 VSS.n207 VSS.n206 5.2005
R3165 VSS.n208 VSS.n207 5.2005
R3166 VSS.n203 VSS.n202 5.2005
R3167 VSS.n209 VSS.n203 5.2005
R3168 VSS.n212 VSS.n211 5.2005
R3169 VSS.n211 VSS.n210 5.2005
R3170 VSS.n213 VSS.n201 5.2005
R3171 VSS.n201 VSS.n200 5.2005
R3172 VSS.n216 VSS.n215 5.2005
R3173 VSS.n217 VSS.n216 5.2005
R3174 VSS.n214 VSS.n199 5.2005
R3175 VSS.n218 VSS.n199 5.2005
R3176 VSS.n220 VSS.n198 5.2005
R3177 VSS.n220 VSS.n219 5.2005
R3178 VSS.n222 VSS.n221 5.2005
R3179 VSS.n221 VSS.n188 5.2005
R3180 VSS.n2818 VSS.n2817 5.2005
R3181 VSS.n2819 VSS.n2818 5.2005
R3182 VSS.n2816 VSS.n197 5.2005
R3183 VSS.n197 VSS.n195 5.2005
R3184 VSS.n2815 VSS.n2814 5.2005
R3185 VSS.n2814 VSS.n2813 5.2005
R3186 VSS.n225 VSS.n224 5.2005
R3187 VSS.n2812 VSS.n225 5.2005
R3188 VSS.n2810 VSS.n2809 5.2005
R3189 VSS.n2811 VSS.n2810 5.2005
R3190 VSS.n2808 VSS.n227 5.2005
R3191 VSS.n227 VSS.n226 5.2005
R3192 VSS.n2807 VSS.n2806 5.2005
R3193 VSS.n2806 VSS.n2805 5.2005
R3194 VSS.n229 VSS.n228 5.2005
R3195 VSS.n2804 VSS.n229 5.2005
R3196 VSS.n2802 VSS.n2801 5.2005
R3197 VSS.n2803 VSS.n2802 5.2005
R3198 VSS.n2800 VSS.n231 5.2005
R3199 VSS.n231 VSS.n230 5.2005
R3200 VSS.n2799 VSS.n2798 5.2005
R3201 VSS.n2798 VSS.n2797 5.2005
R3202 VSS.n233 VSS.n232 5.2005
R3203 VSS.n2796 VSS.n233 5.2005
R3204 VSS.n2794 VSS.n2793 5.2005
R3205 VSS.n2795 VSS.n2794 5.2005
R3206 VSS.n2792 VSS.n235 5.2005
R3207 VSS.n235 VSS.n234 5.2005
R3208 VSS.n2791 VSS.n2790 5.2005
R3209 VSS.n2790 VSS.n2789 5.2005
R3210 VSS.n237 VSS.n236 5.2005
R3211 VSS.n2788 VSS.n237 5.2005
R3212 VSS.n2786 VSS.n2785 5.2005
R3213 VSS.n2787 VSS.n2786 5.2005
R3214 VSS.n2784 VSS.n238 5.2005
R3215 VSS.n241 VSS.n238 5.2005
R3216 VSS.n2783 VSS.n2782 5.2005
R3217 VSS.n2782 VSS.n2781 5.2005
R3218 VSS.n2778 VSS.n2777 5.2005
R3219 VSS.n2779 VSS.n2778 5.2005
R3220 VSS.n2776 VSS.n2774 5.2005
R3221 VSS.n2774 VSS.n2773 5.2005
R3222 VSS.n2775 VSS.n163 5.2005
R3223 VSS.n164 VSS.n163 5.2005
R3224 VSS.n3118 VSS.n162 5.2005
R3225 VSS.n3118 VSS.n3117 5.2005
R3226 VSS.n3121 VSS.n3120 5.2005
R3227 VSS.n3122 VSS.n161 5.2005
R3228 VSS.n3124 VSS.n3123 5.2005
R3229 VSS.n3124 VSS.n98 5.2005
R3230 VSS.n3125 VSS.n160 5.2005
R3231 VSS.n3128 VSS.n3127 5.2005
R3232 VSS.n3129 VSS.n159 5.2005
R3233 VSS.n159 VSS.n98 5.2005
R3234 VSS.n3131 VSS.n3130 5.2005
R3235 VSS.n3133 VSS.n158 5.2005
R3236 VSS.n3134 VSS.n157 5.2005
R3237 VSS.n3134 VSS.n100 5.2005
R3238 VSS.n3137 VSS.n3136 5.2005
R3239 VSS.n3138 VSS.n156 5.2005
R3240 VSS.n3140 VSS.n3139 5.2005
R3241 VSS.n3142 VSS.n155 5.2005
R3242 VSS.n3143 VSS.n154 5.2005
R3243 VSS.n3146 VSS.n3145 5.2005
R3244 VSS.n3149 VSS.n3148 5.2005
R3245 VSS.n3151 VSS.n151 5.2005
R3246 VSS.n3154 VSS.n3153 5.2005
R3247 VSS.n3155 VSS.n150 5.2005
R3248 VSS.n3157 VSS.n3156 5.2005
R3249 VSS.n3159 VSS.n149 5.2005
R3250 VSS.n3162 VSS.n3161 5.2005
R3251 VSS.n3163 VSS.n148 5.2005
R3252 VSS.n3165 VSS.n3164 5.2005
R3253 VSS.n3167 VSS.n147 5.2005
R3254 VSS.n3170 VSS.n3169 5.2005
R3255 VSS.n3171 VSS.n146 5.2005
R3256 VSS.n3173 VSS.n3172 5.2005
R3257 VSS.n3175 VSS.n145 5.2005
R3258 VSS.n3178 VSS.n3177 5.2005
R3259 VSS.n3179 VSS.n144 5.2005
R3260 VSS.n3181 VSS.n3180 5.2005
R3261 VSS.n3183 VSS.n143 5.2005
R3262 VSS.n3185 VSS.n3184 5.2005
R3263 VSS.n3184 VSS.n100 5.2005
R3264 VSS.n3242 VSS.n3241 5.15774
R3265 VSS.n2448 VSS.n2446 4.74734
R3266 VSS.n2635 VSS.n2633 4.51084
R3267 VSS.n3117 VSS.n3116 4.50813
R3268 VSS.n1397 VSS.n1372 4.5005
R3269 VSS.n1408 VSS.n1372 4.5005
R3270 VSS.n1386 VSS.n1372 4.5005
R3271 VSS.n1411 VSS.n1372 4.5005
R3272 VSS.n1384 VSS.n1372 4.5005
R3273 VSS.n1414 VSS.n1372 4.5005
R3274 VSS.n1383 VSS.n1372 4.5005
R3275 VSS.n1416 VSS.n1372 4.5005
R3276 VSS.n1386 VSS.n1286 4.5005
R3277 VSS.n1411 VSS.n1286 4.5005
R3278 VSS.n1384 VSS.n1286 4.5005
R3279 VSS.n1414 VSS.n1286 4.5005
R3280 VSS.n1383 VSS.n1286 4.5005
R3281 VSS.n1416 VSS.n1286 4.5005
R3282 VSS.n1418 VSS.n1286 4.5005
R3283 VSS.n1386 VSS.n1363 4.5005
R3284 VSS.n1411 VSS.n1363 4.5005
R3285 VSS.n1384 VSS.n1363 4.5005
R3286 VSS.n1414 VSS.n1363 4.5005
R3287 VSS.n1383 VSS.n1363 4.5005
R3288 VSS.n1416 VSS.n1363 4.5005
R3289 VSS.n1418 VSS.n1363 4.5005
R3290 VSS.n1386 VSS.n1375 4.5005
R3291 VSS.n1411 VSS.n1375 4.5005
R3292 VSS.n1384 VSS.n1375 4.5005
R3293 VSS.n1414 VSS.n1375 4.5005
R3294 VSS.n1383 VSS.n1375 4.5005
R3295 VSS.n1416 VSS.n1375 4.5005
R3296 VSS.n1418 VSS.n1375 4.5005
R3297 VSS.n1386 VSS.n1362 4.5005
R3298 VSS.n1411 VSS.n1362 4.5005
R3299 VSS.n1384 VSS.n1362 4.5005
R3300 VSS.n1414 VSS.n1362 4.5005
R3301 VSS.n1383 VSS.n1362 4.5005
R3302 VSS.n1416 VSS.n1362 4.5005
R3303 VSS.n1418 VSS.n1362 4.5005
R3304 VSS.n1386 VSS.n1376 4.5005
R3305 VSS.n1411 VSS.n1376 4.5005
R3306 VSS.n1384 VSS.n1376 4.5005
R3307 VSS.n1414 VSS.n1376 4.5005
R3308 VSS.n1383 VSS.n1376 4.5005
R3309 VSS.n1416 VSS.n1376 4.5005
R3310 VSS.n1418 VSS.n1376 4.5005
R3311 VSS.n1386 VSS.n1361 4.5005
R3312 VSS.n1411 VSS.n1361 4.5005
R3313 VSS.n1384 VSS.n1361 4.5005
R3314 VSS.n1414 VSS.n1361 4.5005
R3315 VSS.n1383 VSS.n1361 4.5005
R3316 VSS.n1416 VSS.n1361 4.5005
R3317 VSS.n1418 VSS.n1361 4.5005
R3318 VSS.n1386 VSS.n1377 4.5005
R3319 VSS.n1411 VSS.n1377 4.5005
R3320 VSS.n1384 VSS.n1377 4.5005
R3321 VSS.n1414 VSS.n1377 4.5005
R3322 VSS.n1383 VSS.n1377 4.5005
R3323 VSS.n1416 VSS.n1377 4.5005
R3324 VSS.n1418 VSS.n1377 4.5005
R3325 VSS.n1386 VSS.n1360 4.5005
R3326 VSS.n1411 VSS.n1360 4.5005
R3327 VSS.n1384 VSS.n1360 4.5005
R3328 VSS.n1414 VSS.n1360 4.5005
R3329 VSS.n1383 VSS.n1360 4.5005
R3330 VSS.n1416 VSS.n1360 4.5005
R3331 VSS.n1418 VSS.n1360 4.5005
R3332 VSS.n1386 VSS.n1378 4.5005
R3333 VSS.n1411 VSS.n1378 4.5005
R3334 VSS.n1384 VSS.n1378 4.5005
R3335 VSS.n1414 VSS.n1378 4.5005
R3336 VSS.n1383 VSS.n1378 4.5005
R3337 VSS.n1416 VSS.n1378 4.5005
R3338 VSS.n1418 VSS.n1378 4.5005
R3339 VSS.n1386 VSS.n1359 4.5005
R3340 VSS.n1411 VSS.n1359 4.5005
R3341 VSS.n1384 VSS.n1359 4.5005
R3342 VSS.n1414 VSS.n1359 4.5005
R3343 VSS.n1383 VSS.n1359 4.5005
R3344 VSS.n1416 VSS.n1359 4.5005
R3345 VSS.n1418 VSS.n1359 4.5005
R3346 VSS.n1386 VSS.n1379 4.5005
R3347 VSS.n1411 VSS.n1379 4.5005
R3348 VSS.n1384 VSS.n1379 4.5005
R3349 VSS.n1414 VSS.n1379 4.5005
R3350 VSS.n1383 VSS.n1379 4.5005
R3351 VSS.n1416 VSS.n1379 4.5005
R3352 VSS.n1418 VSS.n1379 4.5005
R3353 VSS.n1386 VSS.n1358 4.5005
R3354 VSS.n1411 VSS.n1358 4.5005
R3355 VSS.n1384 VSS.n1358 4.5005
R3356 VSS.n1414 VSS.n1358 4.5005
R3357 VSS.n1383 VSS.n1358 4.5005
R3358 VSS.n1416 VSS.n1358 4.5005
R3359 VSS.n1418 VSS.n1358 4.5005
R3360 VSS.n1386 VSS.n1380 4.5005
R3361 VSS.n1411 VSS.n1380 4.5005
R3362 VSS.n1384 VSS.n1380 4.5005
R3363 VSS.n1414 VSS.n1380 4.5005
R3364 VSS.n1383 VSS.n1380 4.5005
R3365 VSS.n1416 VSS.n1380 4.5005
R3366 VSS.n1418 VSS.n1380 4.5005
R3367 VSS.n1386 VSS.n1357 4.5005
R3368 VSS.n1411 VSS.n1357 4.5005
R3369 VSS.n1384 VSS.n1357 4.5005
R3370 VSS.n1414 VSS.n1357 4.5005
R3371 VSS.n1383 VSS.n1357 4.5005
R3372 VSS.n1416 VSS.n1357 4.5005
R3373 VSS.n1418 VSS.n1357 4.5005
R3374 VSS.n1386 VSS.n1381 4.5005
R3375 VSS.n1411 VSS.n1381 4.5005
R3376 VSS.n1384 VSS.n1381 4.5005
R3377 VSS.n1414 VSS.n1381 4.5005
R3378 VSS.n1383 VSS.n1381 4.5005
R3379 VSS.n1416 VSS.n1381 4.5005
R3380 VSS.n1418 VSS.n1381 4.5005
R3381 VSS.n1418 VSS.n1356 4.5005
R3382 VSS.n1417 VSS.n1408 4.5005
R3383 VSS.n1417 VSS.n1386 4.5005
R3384 VSS.n1417 VSS.n1411 4.5005
R3385 VSS.n1417 VSS.n1384 4.5005
R3386 VSS.n1417 VSS.n1414 4.5005
R3387 VSS.n1417 VSS.n1383 4.5005
R3388 VSS.n1417 VSS.n1416 4.5005
R3389 VSS.n1418 VSS.n1417 4.5005
R3390 VSS.n1408 VSS.n1268 4.5005
R3391 VSS.n1386 VSS.n1268 4.5005
R3392 VSS.n1411 VSS.n1268 4.5005
R3393 VSS.n1384 VSS.n1268 4.5005
R3394 VSS.n1414 VSS.n1268 4.5005
R3395 VSS.n1383 VSS.n1268 4.5005
R3396 VSS.n1416 VSS.n1268 4.5005
R3397 VSS.n1418 VSS.n1268 4.5005
R3398 VSS.n1408 VSS.n1291 4.5005
R3399 VSS.n1411 VSS.n1291 4.5005
R3400 VSS.n1384 VSS.n1291 4.5005
R3401 VSS.n1414 VSS.n1291 4.5005
R3402 VSS.n1383 VSS.n1291 4.5005
R3403 VSS.n1416 VSS.n1291 4.5005
R3404 VSS.n1418 VSS.n1291 4.5005
R3405 VSS.n1411 VSS.n1374 4.5005
R3406 VSS.n1384 VSS.n1374 4.5005
R3407 VSS.n1414 VSS.n1374 4.5005
R3408 VSS.n1383 VSS.n1374 4.5005
R3409 VSS.n1416 VSS.n1374 4.5005
R3410 VSS.n1418 VSS.n1374 4.5005
R3411 VSS.n1418 VSS.n1372 4.5005
R3412 VSS.n1371 VSS.n1292 4.5005
R3413 VSS.n1454 VSS.n1246 4.5005
R3414 VSS.n1454 VSS.n1288 4.5005
R3415 VSS.n1454 VSS.n1292 4.5005
R3416 VSS.n1454 VSS.n1453 4.5005
R3417 VSS.n1295 VSS.n1246 4.5005
R3418 VSS.n1369 VSS.n1295 4.5005
R3419 VSS.n1367 VSS.n1295 4.5005
R3420 VSS.n1366 VSS.n1295 4.5005
R3421 VSS.n1364 VSS.n1295 4.5005
R3422 VSS.n1295 VSS.n1288 4.5005
R3423 VSS.n1295 VSS.n1292 4.5005
R3424 VSS.n1453 VSS.n1295 4.5005
R3425 VSS.n1465 VSS.n1464 4.5005
R3426 VSS.n1466 VSS.n1465 4.5005
R3427 VSS.n1468 VSS.n1255 4.5005
R3428 VSS.n1464 VSS.n1255 4.5005
R3429 VSS.n1466 VSS.n1255 4.5005
R3430 VSS.n1468 VSS.n1257 4.5005
R3431 VSS.n1267 VSS.n1257 4.5005
R3432 VSS.n1270 VSS.n1257 4.5005
R3433 VSS.n1266 VSS.n1257 4.5005
R3434 VSS.n1272 VSS.n1257 4.5005
R3435 VSS.n1464 VSS.n1257 4.5005
R3436 VSS.n1466 VSS.n1257 4.5005
R3437 VSS.n1468 VSS.n1254 4.5005
R3438 VSS.n1267 VSS.n1254 4.5005
R3439 VSS.n1270 VSS.n1254 4.5005
R3440 VSS.n1266 VSS.n1254 4.5005
R3441 VSS.n1272 VSS.n1254 4.5005
R3442 VSS.n1464 VSS.n1254 4.5005
R3443 VSS.n1466 VSS.n1254 4.5005
R3444 VSS.n1468 VSS.n1258 4.5005
R3445 VSS.n1267 VSS.n1258 4.5005
R3446 VSS.n1270 VSS.n1258 4.5005
R3447 VSS.n1266 VSS.n1258 4.5005
R3448 VSS.n1272 VSS.n1258 4.5005
R3449 VSS.n1464 VSS.n1258 4.5005
R3450 VSS.n1466 VSS.n1258 4.5005
R3451 VSS.n1468 VSS.n1253 4.5005
R3452 VSS.n1267 VSS.n1253 4.5005
R3453 VSS.n1270 VSS.n1253 4.5005
R3454 VSS.n1266 VSS.n1253 4.5005
R3455 VSS.n1272 VSS.n1253 4.5005
R3456 VSS.n1464 VSS.n1253 4.5005
R3457 VSS.n1466 VSS.n1253 4.5005
R3458 VSS.n1468 VSS.n1259 4.5005
R3459 VSS.n1267 VSS.n1259 4.5005
R3460 VSS.n1270 VSS.n1259 4.5005
R3461 VSS.n1266 VSS.n1259 4.5005
R3462 VSS.n1272 VSS.n1259 4.5005
R3463 VSS.n1464 VSS.n1259 4.5005
R3464 VSS.n1466 VSS.n1259 4.5005
R3465 VSS.n1468 VSS.n1252 4.5005
R3466 VSS.n1267 VSS.n1252 4.5005
R3467 VSS.n1270 VSS.n1252 4.5005
R3468 VSS.n1266 VSS.n1252 4.5005
R3469 VSS.n1272 VSS.n1252 4.5005
R3470 VSS.n1464 VSS.n1252 4.5005
R3471 VSS.n1466 VSS.n1252 4.5005
R3472 VSS.n1468 VSS.n1260 4.5005
R3473 VSS.n1267 VSS.n1260 4.5005
R3474 VSS.n1270 VSS.n1260 4.5005
R3475 VSS.n1266 VSS.n1260 4.5005
R3476 VSS.n1272 VSS.n1260 4.5005
R3477 VSS.n1464 VSS.n1260 4.5005
R3478 VSS.n1466 VSS.n1260 4.5005
R3479 VSS.n1468 VSS.n1251 4.5005
R3480 VSS.n1267 VSS.n1251 4.5005
R3481 VSS.n1270 VSS.n1251 4.5005
R3482 VSS.n1266 VSS.n1251 4.5005
R3483 VSS.n1272 VSS.n1251 4.5005
R3484 VSS.n1464 VSS.n1251 4.5005
R3485 VSS.n1466 VSS.n1251 4.5005
R3486 VSS.n1468 VSS.n1261 4.5005
R3487 VSS.n1267 VSS.n1261 4.5005
R3488 VSS.n1270 VSS.n1261 4.5005
R3489 VSS.n1266 VSS.n1261 4.5005
R3490 VSS.n1272 VSS.n1261 4.5005
R3491 VSS.n1464 VSS.n1261 4.5005
R3492 VSS.n1466 VSS.n1261 4.5005
R3493 VSS.n1468 VSS.n1250 4.5005
R3494 VSS.n1267 VSS.n1250 4.5005
R3495 VSS.n1270 VSS.n1250 4.5005
R3496 VSS.n1266 VSS.n1250 4.5005
R3497 VSS.n1272 VSS.n1250 4.5005
R3498 VSS.n1464 VSS.n1250 4.5005
R3499 VSS.n1466 VSS.n1250 4.5005
R3500 VSS.n1468 VSS.n1262 4.5005
R3501 VSS.n1267 VSS.n1262 4.5005
R3502 VSS.n1270 VSS.n1262 4.5005
R3503 VSS.n1266 VSS.n1262 4.5005
R3504 VSS.n1272 VSS.n1262 4.5005
R3505 VSS.n1464 VSS.n1262 4.5005
R3506 VSS.n1466 VSS.n1262 4.5005
R3507 VSS.n1468 VSS.n1249 4.5005
R3508 VSS.n1267 VSS.n1249 4.5005
R3509 VSS.n1270 VSS.n1249 4.5005
R3510 VSS.n1266 VSS.n1249 4.5005
R3511 VSS.n1272 VSS.n1249 4.5005
R3512 VSS.n1464 VSS.n1249 4.5005
R3513 VSS.n1466 VSS.n1249 4.5005
R3514 VSS.n1468 VSS.n1263 4.5005
R3515 VSS.n1267 VSS.n1263 4.5005
R3516 VSS.n1270 VSS.n1263 4.5005
R3517 VSS.n1266 VSS.n1263 4.5005
R3518 VSS.n1272 VSS.n1263 4.5005
R3519 VSS.n1464 VSS.n1263 4.5005
R3520 VSS.n1466 VSS.n1263 4.5005
R3521 VSS.n1468 VSS.n1248 4.5005
R3522 VSS.n1267 VSS.n1248 4.5005
R3523 VSS.n1270 VSS.n1248 4.5005
R3524 VSS.n1266 VSS.n1248 4.5005
R3525 VSS.n1272 VSS.n1248 4.5005
R3526 VSS.n1464 VSS.n1248 4.5005
R3527 VSS.n1466 VSS.n1248 4.5005
R3528 VSS.n1468 VSS.n1264 4.5005
R3529 VSS.n1267 VSS.n1264 4.5005
R3530 VSS.n1270 VSS.n1264 4.5005
R3531 VSS.n1266 VSS.n1264 4.5005
R3532 VSS.n1272 VSS.n1264 4.5005
R3533 VSS.n1464 VSS.n1264 4.5005
R3534 VSS.n1466 VSS.n1264 4.5005
R3535 VSS.n1468 VSS.n1247 4.5005
R3536 VSS.n1267 VSS.n1247 4.5005
R3537 VSS.n1270 VSS.n1247 4.5005
R3538 VSS.n1266 VSS.n1247 4.5005
R3539 VSS.n1272 VSS.n1247 4.5005
R3540 VSS.n1464 VSS.n1247 4.5005
R3541 VSS.n1466 VSS.n1247 4.5005
R3542 VSS.n1468 VSS.n1467 4.5005
R3543 VSS.n1467 VSS.n1267 4.5005
R3544 VSS.n1467 VSS.n1270 4.5005
R3545 VSS.n1467 VSS.n1266 4.5005
R3546 VSS.n1467 VSS.n1272 4.5005
R3547 VSS.n1467 VSS.n1466 4.5005
R3548 VSS.n1451 VSS.n1450 4.5005
R3549 VSS.n1449 VSS.n1299 4.5005
R3550 VSS.n1448 VSS.n1447 4.5005
R3551 VSS.n1446 VSS.n1300 4.5005
R3552 VSS.n1445 VSS.n1444 4.5005
R3553 VSS.n1443 VSS.n1307 4.5005
R3554 VSS.n1442 VSS.n1441 4.5005
R3555 VSS.n1440 VSS.n1308 4.5005
R3556 VSS.n1439 VSS.n1438 4.5005
R3557 VSS.n1437 VSS.n1316 4.5005
R3558 VSS.n1436 VSS.n1435 4.5005
R3559 VSS.n1434 VSS.n1317 4.5005
R3560 VSS.n1433 VSS.n1432 4.5005
R3561 VSS.n1431 VSS.n1325 4.5005
R3562 VSS.n1430 VSS.n1429 4.5005
R3563 VSS.n1428 VSS.n1326 4.5005
R3564 VSS.n1427 VSS.n1426 4.5005
R3565 VSS.n1425 VSS.n1424 4.5005
R3566 VSS.n1421 VSS.n103 4.5005
R3567 VSS.n3233 VSS.n3228 4.43655
R3568 VSS.n1809 VSS.n900 4.43088
R3569 VSS.n1807 VSS.n1806 4.43088
R3570 VSS.n1804 VSS.n903 4.43088
R3571 VSS.n1800 VSS.n1798 4.43088
R3572 VSS.n1794 VSS.n1793 4.43088
R3573 VSS.n1791 VSS.n909 4.43088
R3574 VSS.n1787 VSS.n909 4.43088
R3575 VSS.n920 VSS.n911 4.43088
R3576 VSS.n1591 VSS.n1589 4.43088
R3577 VSS.n1591 VSS.n1587 4.43088
R3578 VSS.n1595 VSS.n1587 4.43088
R3579 VSS.n1595 VSS.n1585 4.43088
R3580 VSS.n1600 VSS.n1585 4.43088
R3581 VSS.n1600 VSS.n1583 4.43088
R3582 VSS.n1604 VSS.n1583 4.43088
R3583 VSS.n1605 VSS.n1604 4.43088
R3584 VSS.n1605 VSS.n1582 4.43088
R3585 VSS.n1609 VSS.n1582 4.43088
R3586 VSS.n1609 VSS.n1580 4.43088
R3587 VSS.n1613 VSS.n1580 4.43088
R3588 VSS.n1613 VSS.n1577 4.43088
R3589 VSS.n1624 VSS.n1577 4.43088
R3590 VSS.n1624 VSS.n1578 4.43088
R3591 VSS.n1620 VSS.n1619 4.43088
R3592 VSS.n2635 VSS.n2634 4.38259
R3593 VSS.t83 VSS.t144 4.27307
R3594 VSS.n1179 VSS.n1178 4.13154
R3595 VSS.n1517 VSS.n994 4.12546
R3596 VSS.n1520 VSS.n994 4.12546
R3597 VSS.n142 VSS.n109 4.11885
R3598 VSS.n944 VSS.t299 4.0955
R3599 VSS.n1683 VSS.t198 4.0955
R3600 VSS.n1682 VSS.t151 4.0955
R3601 VSS.n1888 VSS.n1887 4.05793
R3602 VSS.n2060 VSS.n2059 4.05793
R3603 VSS.n2165 VSS.n2164 4.05793
R3604 VSS.n2337 VSS.n2336 4.05793
R3605 VSS.n470 VSS.n191 4.05793
R3606 VSS.n941 VSS.t32 4.04494
R3607 VSS.n941 VSS.t234 4.04494
R3608 VSS.n1687 VSS.t291 4.04494
R3609 VSS.n1687 VSS.t205 4.04494
R3610 VSS.n1686 VSS.t302 4.04494
R3611 VSS.n1686 VSS.t200 4.04494
R3612 VSS.n930 VSS.t232 4.04494
R3613 VSS.n930 VSS.t237 4.04494
R3614 VSS.n1727 VSS.n1726 3.89923
R3615 VSS.n1796 VSS.n906 3.8975
R3616 VSS.n1698 VSS.t96 3.8098
R3617 VSS.n1698 VSS.t100 3.8098
R3618 VSS.n1699 VSS.t88 3.8098
R3619 VSS.n1699 VSS.t98 3.8098
R3620 VSS.n1700 VSS.t102 3.8098
R3621 VSS.n1700 VSS.t90 3.8098
R3622 VSS.n1545 VSS.n1001 3.80605
R3623 VSS.n1541 VSS.n1000 3.80605
R3624 VSS.n1537 VSS.n999 3.80605
R3625 VSS.n1533 VSS.n998 3.80605
R3626 VSS.n1529 VSS.n997 3.80605
R3627 VSS.n1525 VSS.n996 3.80605
R3628 VSS.n1521 VSS.n995 3.80605
R3629 VSS.n1524 VSS.n995 3.80605
R3630 VSS.n1528 VSS.n996 3.80605
R3631 VSS.n1532 VSS.n997 3.80605
R3632 VSS.n1536 VSS.n998 3.80605
R3633 VSS.n1540 VSS.n999 3.80605
R3634 VSS.n1544 VSS.n1000 3.80605
R3635 VSS.n1003 VSS.n1001 3.80605
R3636 VSS.n1059 VSS.n1058 3.79267
R3637 VSS.n1054 VSS.n1024 3.79267
R3638 VSS.n1052 VSS.n1051 3.79267
R3639 VSS.n1047 VSS.n1027 3.79267
R3640 VSS.n1045 VSS.n1044 3.79267
R3641 VSS.n1040 VSS.n1030 3.79267
R3642 VSS.n1038 VSS.n1037 3.79267
R3643 VSS.n1033 VSS.n1032 3.79267
R3644 VSS.n1197 VSS.n1196 3.79267
R3645 VSS.n1126 VSS.n1087 3.79267
R3646 VSS.n1130 VSS.n1088 3.79267
R3647 VSS.n1134 VSS.n1089 3.79267
R3648 VSS.n1138 VSS.n1090 3.79267
R3649 VSS.n1142 VSS.n1091 3.79267
R3650 VSS.n1146 VSS.n1092 3.79267
R3651 VSS.n1150 VSS.n1093 3.79267
R3652 VSS.n1197 VSS.n1096 3.79267
R3653 VSS.n1129 VSS.n1087 3.79267
R3654 VSS.n1133 VSS.n1088 3.79267
R3655 VSS.n1137 VSS.n1089 3.79267
R3656 VSS.n1141 VSS.n1090 3.79267
R3657 VSS.n1145 VSS.n1091 3.79267
R3658 VSS.n1149 VSS.n1092 3.79267
R3659 VSS.n1155 VSS.n1093 3.79267
R3660 VSS.n1032 VSS.n1031 3.79267
R3661 VSS.n1039 VSS.n1038 3.79267
R3662 VSS.n1030 VSS.n1028 3.79267
R3663 VSS.n1046 VSS.n1045 3.79267
R3664 VSS.n1027 VSS.n1025 3.79267
R3665 VSS.n1053 VSS.n1052 3.79267
R3666 VSS.n1024 VSS.n1022 3.79267
R3667 VSS.n1060 VSS.n1059 3.79267
R3668 VSS.n3194 VSS.n107 3.73488
R3669 VSS.n1847 VSS.n23 3.71266
R3670 VSS.n45 VSS.n40 3.71266
R3671 VSS.n67 VSS.n62 3.71266
R3672 VSS.n89 VSS.n84 3.71266
R3673 VSS.n2821 VSS.n2820 3.71266
R3674 VSS.t284 VSS.t233 3.71055
R3675 VSS.n3199 VSS.n127 3.69405
R3676 VSS.n3198 VSS.n3189 3.69405
R3677 VSS.n3187 VSS.n3186 3.69405
R3678 VSS.n1187 VSS.n1186 3.64321
R3679 VSS.n1186 VSS.n1185 3.64321
R3680 VSS.n929 VSS.t178 3.6005
R3681 VSS.n929 VSS.t174 3.6005
R3682 VSS.n2748 VSS.n260 3.59261
R3683 VSS.n2487 VSS.n478 3.59261
R3684 VSS.n2341 VSS.n535 3.59261
R3685 VSS.n2103 VSS.n696 3.59261
R3686 VSS.n2064 VSS.n715 3.59261
R3687 VSS.n350 VSS.n349 3.59261
R3688 VSS.n1877 VSS.n1876 3.59261
R3689 VSS.n247 VSS.n242 3.32459
R3690 VSS.n2772 VSS.n2771 3.32459
R3691 VSS.n2766 VSS.n2765 3.32459
R3692 VSS.n2763 VSS.n2762 3.32459
R3693 VSS.n2758 VSS.n255 3.32459
R3694 VSS.n2756 VSS.n2755 3.32459
R3695 VSS.n2751 VSS.n258 3.32459
R3696 VSS.n2749 VSS.n2748 3.32459
R3697 VSS.n487 VSS.n189 3.32459
R3698 VSS.n491 VSS.n190 3.32459
R3699 VSS.n493 VSS.n482 3.32459
R3700 VSS.n500 VSS.n499 3.32459
R3701 VSS.n501 VSS.n480 3.32459
R3702 VSS.n508 VSS.n507 3.32459
R3703 VSS.n511 VSS.n476 3.32459
R3704 VSS.n2488 VSS.n2487 3.32459
R3705 VSS.n557 VSS.n556 3.32459
R3706 VSS.n558 VSS.n552 3.32459
R3707 VSS.n571 VSS.n551 3.32459
R3708 VSS.n567 VSS.n550 3.32459
R3709 VSS.n563 VSS.n549 3.32459
R3710 VSS.n578 VSS.n577 3.32459
R3711 VSS.n582 VSS.n542 3.32459
R3712 VSS.n543 VSS.n535 3.32459
R3713 VSS.n1880 VSS.n831 3.32459
R3714 VSS.n1885 VSS.n1884 3.32459
R3715 VSS.n813 VSS.n812 3.32459
R3716 VSS.n1922 VSS.n1921 3.32459
R3717 VSS.n768 VSS.n721 3.32459
R3718 VSS.n724 VSS.n722 3.32459
R3719 VSS.n2029 VSS.n2028 3.32459
R3720 VSS.n2026 VSS.n2025 3.32459
R3721 VSS.n2162 VSS.n2161 3.32459
R3722 VSS.n2157 VSS.n652 3.32459
R3723 VSS.n634 VSS.n633 3.32459
R3724 VSS.n2199 VSS.n2198 3.32459
R3725 VSS.n589 VSS.n540 3.32459
R3726 VSS.n545 VSS.n541 3.32459
R3727 VSS.n2306 VSS.n2305 3.32459
R3728 VSS.n2303 VSS.n2302 3.32459
R3729 VSS.n514 VSS.n475 3.32459
R3730 VSS.n2491 VSS.n2490 3.32459
R3731 VSS.n2520 VSS.n454 3.32459
R3732 VSS.n456 VSS.n455 3.32459
R3733 VSS.n1922 VSS.n1920 3.32459
R3734 VSS.n1916 VSS.n812 3.32459
R3735 VSS.n2027 VSS.n2026 3.32459
R3736 VSS.n2030 VSS.n2029 3.32459
R3737 VSS.n2199 VSS.n2197 3.32459
R3738 VSS.n2193 VSS.n633 3.32459
R3739 VSS.n2304 VSS.n2303 3.32459
R3740 VSS.n2307 VSS.n2306 3.32459
R3741 VSS.n2519 VSS.n456 3.32459
R3742 VSS.n459 VSS.n454 3.32459
R3743 VSS.n583 VSS.n543 3.32459
R3744 VSS.n579 VSS.n542 3.32459
R3745 VSS.n2488 VSS.n477 3.32459
R3746 VSS.n509 VSS.n476 3.32459
R3747 VSS.n2750 VSS.n2749 3.32459
R3748 VSS.n258 VSS.n256 3.32459
R3749 VSS.n1885 VSS.n832 3.32459
R3750 VSS.n1878 VSS.n831 3.32459
R3751 VSS.n769 VSS.n722 3.32459
R3752 VSS.n721 VSS.n714 3.32459
R3753 VSS.n654 VSS.n652 3.32459
R3754 VSS.n2162 VSS.n653 3.32459
R3755 VSS.n590 VSS.n541 3.32459
R3756 VSS.n540 VSS.n536 3.32459
R3757 VSS.n2490 VSS.n473 3.32459
R3758 VSS.n516 VSS.n475 3.32459
R3759 VSS.n665 VSS.n664 3.32459
R3760 VSS.n666 VSS.n660 3.32459
R3761 VSS.n679 VSS.n659 3.32459
R3762 VSS.n675 VSS.n658 3.32459
R3763 VSS.n671 VSS.n657 3.32459
R3764 VSS.n686 VSS.n685 3.32459
R3765 VSS.n687 VSS.n650 3.32459
R3766 VSS.n691 VSS.n651 3.32459
R3767 VSS.n696 VSS.n651 3.32459
R3768 VSS.n690 VSS.n650 3.32459
R3769 VSS.n685 VSS.n656 3.32459
R3770 VSS.n674 VSS.n657 3.32459
R3771 VSS.n678 VSS.n658 3.32459
R3772 VSS.n661 VSS.n659 3.32459
R3773 VSS.n577 VSS.n548 3.32459
R3774 VSS.n566 VSS.n549 3.32459
R3775 VSS.n570 VSS.n550 3.32459
R3776 VSS.n553 VSS.n551 3.32459
R3777 VSS.n507 VSS.n506 3.32459
R3778 VSS.n502 VSS.n501 3.32459
R3779 VSS.n499 VSS.n498 3.32459
R3780 VSS.n494 VSS.n493 3.32459
R3781 VSS.n2757 VSS.n2756 3.32459
R3782 VSS.n255 VSS.n253 3.32459
R3783 VSS.n2764 VSS.n2763 3.32459
R3784 VSS.n2767 VSS.n2766 3.32459
R3785 VSS.n2405 VSS.n2404 3.32459
R3786 VSS.n2406 VSS.n2400 3.32459
R3787 VSS.n2577 VSS.n426 3.32459
R3788 VSS.n2580 VSS.n2579 3.32459
R3789 VSS.n2579 VSS.n2578 3.32459
R3790 VSS.n2574 VSS.n426 3.32459
R3791 VSS.n2407 VSS.n2406 3.32459
R3792 VSS.n2404 VSS.n2403 3.32459
R3793 VSS.n736 VSS.n735 3.32459
R3794 VSS.n737 VSS.n731 3.32459
R3795 VSS.n750 VSS.n730 3.32459
R3796 VSS.n746 VSS.n729 3.32459
R3797 VSS.n742 VSS.n728 3.32459
R3798 VSS.n757 VSS.n756 3.32459
R3799 VSS.n761 VSS.n719 3.32459
R3800 VSS.n720 VSS.n715 3.32459
R3801 VSS.n762 VSS.n720 3.32459
R3802 VSS.n758 VSS.n719 3.32459
R3803 VSS.n756 VSS.n727 3.32459
R3804 VSS.n745 VSS.n728 3.32459
R3805 VSS.n749 VSS.n729 3.32459
R3806 VSS.n732 VSS.n730 3.32459
R3807 VSS.n3120 VSS.n3119 3.32459
R3808 VSS.n3126 VSS.n3125 3.32459
R3809 VSS.n3132 VSS.n3131 3.32459
R3810 VSS.n3136 VSS.n3135 3.32459
R3811 VSS.n3141 VSS.n3140 3.32459
R3812 VSS.n3144 VSS.n3143 3.32459
R3813 VSS.n3150 VSS.n3149 3.32459
R3814 VSS.n3153 VSS.n3152 3.32459
R3815 VSS.n3158 VSS.n3157 3.32459
R3816 VSS.n3161 VSS.n3160 3.32459
R3817 VSS.n3166 VSS.n3165 3.32459
R3818 VSS.n3169 VSS.n3168 3.32459
R3819 VSS.n3174 VSS.n3173 3.32459
R3820 VSS.n3177 VSS.n3176 3.32459
R3821 VSS.n3182 VSS.n3181 3.32459
R3822 VSS.n328 VSS.n327 3.32459
R3823 VSS.n334 VSS.n306 3.32459
R3824 VSS.n341 VSS.n340 3.32459
R3825 VSS.n342 VSS.n304 3.32459
R3826 VSS.n349 VSS.n348 3.32459
R3827 VSS.n348 VSS.n347 3.32459
R3828 VSS.n343 VSS.n342 3.32459
R3829 VSS.n340 VSS.n339 3.32459
R3830 VSS.n335 VSS.n334 3.32459
R3831 VSS.n328 VSS.n309 3.32459
R3832 VSS.n365 VSS.n364 3.32459
R3833 VSS.n362 VSS.n361 3.32459
R3834 VSS.n357 VSS.n354 3.32459
R3835 VSS.n355 VSS.n288 3.32459
R3836 VSS.n2638 VSS.n2623 3.32459
R3837 VSS.n2642 VSS.n2624 3.32459
R3838 VSS.n2626 VSS.n2625 3.32459
R3839 VSS.n2649 VSS.n2648 3.32459
R3840 VSS.n2649 VSS.n2647 3.32459
R3841 VSS.n2643 VSS.n2625 3.32459
R3842 VSS.n2639 VSS.n2624 3.32459
R3843 VSS.n2632 VSS.n2623 3.32459
R3844 VSS.n356 VSS.n355 3.32459
R3845 VSS.n354 VSS.n352 3.32459
R3846 VSS.n363 VSS.n362 3.32459
R3847 VSS.n366 VSS.n365 3.32459
R3848 VSS.n2735 VSS.n2734 3.32459
R3849 VSS.n2732 VSS.n2731 3.32459
R3850 VSS.n3215 VSS.n3214 3.32459
R3851 VSS.n3212 VSS.n3211 3.32459
R3852 VSS.n3207 VSS.n140 3.32459
R3853 VSS.n140 VSS.n138 3.32459
R3854 VSS.n3213 VSS.n3212 3.32459
R3855 VSS.n3216 VSS.n3215 3.32459
R3856 VSS.n2733 VSS.n2732 3.32459
R3857 VSS.n2736 VSS.n2735 3.32459
R3858 VSS.n1846 VSS.n1844 3.32459
R3859 VSS.n1848 VSS.n1841 3.32459
R3860 VSS.n1861 VSS.n1840 3.32459
R3861 VSS.n1857 VSS.n1839 3.32459
R3862 VSS.n1853 VSS.n1838 3.32459
R3863 VSS.n1868 VSS.n1867 3.32459
R3864 VSS.n1872 VSS.n829 3.32459
R3865 VSS.n1876 VSS.n830 3.32459
R3866 VSS.n1873 VSS.n830 3.32459
R3867 VSS.n1869 VSS.n829 3.32459
R3868 VSS.n1867 VSS.n888 3.32459
R3869 VSS.n1856 VSS.n1838 3.32459
R3870 VSS.n1860 VSS.n1839 3.32459
R3871 VSS.n1842 VSS.n1840 3.32459
R3872 VSS.n1849 VSS.n1848 3.32459
R3873 VSS.n1846 VSS.n1845 3.32459
R3874 VSS.n738 VSS.n737 3.32459
R3875 VSS.n735 VSS.n734 3.32459
R3876 VSS.n667 VSS.n666 3.32459
R3877 VSS.n664 VSS.n663 3.32459
R3878 VSS.n559 VSS.n558 3.32459
R3879 VSS.n556 VSS.n555 3.32459
R3880 VSS.n488 VSS.n190 3.32459
R3881 VSS.n484 VSS.n189 3.32459
R3882 VSS.n2772 VSS.n243 3.32459
R3883 VSS.n245 VSS.n242 3.32459
R3884 VSS.n3119 VSS.n161 3.32459
R3885 VSS.n3127 VSS.n3126 3.32459
R3886 VSS.n3133 VSS.n3132 3.32459
R3887 VSS.n3135 VSS.n156 3.32459
R3888 VSS.n3142 VSS.n3141 3.32459
R3889 VSS.n3145 VSS.n3144 3.32459
R3890 VSS.n3151 VSS.n3150 3.32459
R3891 VSS.n3152 VSS.n150 3.32459
R3892 VSS.n3159 VSS.n3158 3.32459
R3893 VSS.n3160 VSS.n148 3.32459
R3894 VSS.n3167 VSS.n3166 3.32459
R3895 VSS.n3168 VSS.n146 3.32459
R3896 VSS.n3175 VSS.n3174 3.32459
R3897 VSS.n3176 VSS.n144 3.32459
R3898 VSS.n3183 VSS.n3182 3.32459
R3899 VSS.n3233 VSS.n3232 3.25471
R3900 VSS.n3199 VSS.n114 3.25471
R3901 VSS.n3198 VSS.n3197 3.25471
R3902 VSS.n1837 VSS.n1836 3.18236
R3903 VSS.n3260 VSS.n3259 3.11113
R3904 VSS.n1201 VSS.t59 3.00489
R3905 VSS.n3249 VSS.n116 2.91603
R3906 VSS.n1729 VSS.n917 2.72518
R3907 VSS.n962 VSS.n961 2.66171
R3908 VSS.n1680 VSS.n927 2.66171
R3909 VSS.n3256 VSS.n108 2.60721
R3910 VSS.n1182 VSS.n1108 2.54316
R3911 VSS.n1181 VSS.n1109 2.54316
R3912 VSS.n1115 VSS.n1108 2.54316
R3913 VSS.n1206 VSS.t28 2.5205
R3914 VSS.n1206 VSS.t248 2.5205
R3915 VSS.n3225 VSS.n128 2.4855
R3916 VSS.n1551 VSS.n1550 2.38689
R3917 VSS.n1452 VSS.n1451 2.2505
R3918 VSS.n1299 VSS.n1296 2.2505
R3919 VSS.n1447 VSS.n1301 2.2505
R3920 VSS.n1446 VSS.n1303 2.2505
R3921 VSS.n1445 VSS.n1305 2.2505
R3922 VSS.n1309 VSS.n1307 2.2505
R3923 VSS.n1441 VSS.n1310 2.2505
R3924 VSS.n1440 VSS.n1312 2.2505
R3925 VSS.n1439 VSS.n1314 2.2505
R3926 VSS.n1318 VSS.n1316 2.2505
R3927 VSS.n1435 VSS.n1319 2.2505
R3928 VSS.n1434 VSS.n1321 2.2505
R3929 VSS.n1433 VSS.n1323 2.2505
R3930 VSS.n1327 VSS.n1325 2.2505
R3931 VSS.n1429 VSS.n1328 2.2505
R3932 VSS.n1428 VSS.n1330 2.2505
R3933 VSS.n1427 VSS.n1332 2.2505
R3934 VSS.n1409 VSS.n1356 2.25002
R3935 VSS.n1412 VSS.n1356 2.25002
R3936 VSS.n1415 VSS.n1356 2.25002
R3937 VSS.n1399 VSS.n1382 2.25002
R3938 VSS.n1410 VSS.n1382 2.25002
R3939 VSS.n1413 VSS.n1382 2.25002
R3940 VSS.n1382 VSS.n1355 2.25002
R3941 VSS.n1398 VSS.n1374 2.25002
R3942 VSS.n1465 VSS.n1256 2.24986
R3943 VSS.n1465 VSS.n1285 2.24986
R3944 VSS.n1465 VSS.n1284 2.24986
R3945 VSS.n1269 VSS.n1255 2.24986
R3946 VSS.n1271 VSS.n1255 2.24986
R3947 VSS.n1467 VSS.n1273 2.24986
R3948 VSS.n1397 VSS.n1396 2.24873
R3949 VSS.n1408 VSS.n1407 2.24873
R3950 VSS.n1397 VSS.n1395 2.24873
R3951 VSS.n1408 VSS.n1406 2.24873
R3952 VSS.n1397 VSS.n1394 2.24873
R3953 VSS.n1408 VSS.n1405 2.24873
R3954 VSS.n1397 VSS.n1393 2.24873
R3955 VSS.n1408 VSS.n1404 2.24873
R3956 VSS.n1397 VSS.n1392 2.24873
R3957 VSS.n1408 VSS.n1403 2.24873
R3958 VSS.n1397 VSS.n1391 2.24873
R3959 VSS.n1408 VSS.n1402 2.24873
R3960 VSS.n1397 VSS.n1390 2.24873
R3961 VSS.n1408 VSS.n1401 2.24873
R3962 VSS.n1397 VSS.n1389 2.24873
R3963 VSS.n1408 VSS.n1400 2.24873
R3964 VSS.n1397 VSS.n1387 2.24873
R3965 VSS.n1397 VSS.n1388 2.24873
R3966 VSS.n1386 VSS.n1385 2.24873
R3967 VSS.n1293 VSS.n1287 2.24873
R3968 VSS.n1283 VSS.n1282 2.24873
R3969 VSS.n1463 VSS.n1462 2.24873
R3970 VSS.n1282 VSS.n1274 2.24873
R3971 VSS.n1463 VSS.n1461 2.24873
R3972 VSS.n1282 VSS.n1275 2.24873
R3973 VSS.n1463 VSS.n1460 2.24873
R3974 VSS.n1282 VSS.n1276 2.24873
R3975 VSS.n1463 VSS.n1459 2.24873
R3976 VSS.n1282 VSS.n1277 2.24873
R3977 VSS.n1463 VSS.n1458 2.24873
R3978 VSS.n1282 VSS.n1278 2.24873
R3979 VSS.n1463 VSS.n1457 2.24873
R3980 VSS.n1282 VSS.n1279 2.24873
R3981 VSS.n1463 VSS.n1456 2.24873
R3982 VSS.n1282 VSS.n1280 2.24873
R3983 VSS.n1463 VSS.n1455 2.24873
R3984 VSS.n1282 VSS.n1281 2.24873
R3985 VSS.n1463 VSS.n1265 2.24873
R3986 VSS.n1371 VSS.n1370 2.24231
R3987 VSS.n1371 VSS.n1368 2.24231
R3988 VSS.n1371 VSS.n1365 2.24231
R3989 VSS.n1454 VSS.n1290 2.24231
R3990 VSS.n1454 VSS.n1289 2.24231
R3991 VSS.n1371 VSS.n1294 2.24231
R3992 VSS.n3262 VSS.n3261 2.219
R3993 VSS.n3423 VSS.n8 2.15937
R3994 VSS.n3427 VSS.n5 2.12174
R3995 VSS.n1114 VSS.t39 2.05866
R3996 VSS.n2823 VSS.n104 1.99927
R3997 VSS.n1114 VSS.t37 1.96984
R3998 VSS.n1204 VSS.t104 1.87824
R3999 VSS.n1786 VSS.n1785 1.82428
R4000 VSS.n1785 VSS.n915 1.82428
R4001 VSS.n1785 VSS.n914 1.82428
R4002 VSS.n1785 VSS.n913 1.82428
R4003 VSS.n1676 VSS.n1570 1.82428
R4004 VSS.n1676 VSS.n1569 1.82428
R4005 VSS.n1805 VSS.n891 1.82428
R4006 VSS.n1799 VSS.n891 1.82428
R4007 VSS.n905 VSS.n891 1.82428
R4008 VSS.n1792 VSS.n891 1.82428
R4009 VSS.n1815 VSS.n1814 1.82428
R4010 VSS.n1815 VSS.n899 1.82428
R4011 VSS.n2636 VSS.n2635 1.81881
R4012 VSS.n1796 VSS.n907 1.80163
R4013 VSS.n1245 VSS.n1244 1.7498
R4014 VSS.n922 VSS.n917 1.7062
R4015 VSS.n1228 VSS.t163 1.6385
R4016 VSS.n1228 VSS.t110 1.6385
R4017 VSS.n1230 VSS.t126 1.6385
R4018 VSS.n1230 VSS.t30 1.6385
R4019 VSS.n3231 VSS.n114 1.58024
R4020 VSS.n3232 VSS.n3231 1.58024
R4021 VSS.n3250 VSS.n3249 1.58024
R4022 VSS.n1814 VSS.n1813 1.55443
R4023 VSS.n1807 VSS.n899 1.55443
R4024 VSS.n1806 VSS.n1805 1.55443
R4025 VSS.n1799 VSS.n903 1.55443
R4026 VSS.n1798 VSS.n905 1.55443
R4027 VSS.n1793 VSS.n1792 1.55443
R4028 VSS.n1787 VSS.n1786 1.55443
R4029 VSS.n920 VSS.n915 1.55443
R4030 VSS.n1729 VSS.n914 1.55443
R4031 VSS.n925 VSS.n913 1.55443
R4032 VSS.n1578 VSS.n1570 1.55443
R4033 VSS.n1619 VSS.n1569 1.55443
R4034 VSS.n1786 VSS.n911 1.55443
R4035 VSS.n922 VSS.n915 1.55443
R4036 VSS.n1727 VSS.n914 1.55443
R4037 VSS.n1589 VSS.n913 1.55443
R4038 VSS.n1620 VSS.n1570 1.55443
R4039 VSS.n1616 VSS.n1569 1.55443
R4040 VSS.n1805 VSS.n1804 1.55443
R4041 VSS.n1800 VSS.n1799 1.55443
R4042 VSS.n1794 VSS.n905 1.55443
R4043 VSS.n1792 VSS.n1791 1.55443
R4044 VSS.n1814 VSS.n900 1.55443
R4045 VSS.n1809 VSS.n899 1.55443
R4046 VSS.n1813 VSS.n897 1.55113
R4047 VSS.n1244 VSS.n1005 1.52481
R4048 VSS.t43 VSS.n1346 1.5005
R4049 VSS.n1419 VSS.n1298 1.5005
R4050 VSS.n1337 VSS.n1336 1.5005
R4051 VSS.n1338 VSS.n1302 1.5005
R4052 VSS.n1339 VSS.n1304 1.5005
R4053 VSS.n1340 VSS.n1306 1.5005
R4054 VSS.n1342 VSS.n1341 1.5005
R4055 VSS.n1343 VSS.n1311 1.5005
R4056 VSS.n1344 VSS.n1313 1.5005
R4057 VSS.n1345 VSS.n1315 1.5005
R4058 VSS.n1354 VSS.n1320 1.5005
R4059 VSS.n1353 VSS.n1322 1.5005
R4060 VSS.n1352 VSS.n1324 1.5005
R4061 VSS.n1351 VSS.n1350 1.5005
R4062 VSS.n1349 VSS.n1329 1.5005
R4063 VSS.n1348 VSS.n1331 1.5005
R4064 VSS.n1347 VSS.n1333 1.5005
R4065 VSS.n1423 VSS.n1335 1.5005
R4066 VSS.n1422 VSS.n1420 1.5005
R4067 VSS.n1451 VSS.n1298 1.5005
R4068 VSS.n1336 VSS.n1299 1.5005
R4069 VSS.n1447 VSS.n1302 1.5005
R4070 VSS.n1446 VSS.n1304 1.5005
R4071 VSS.n1445 VSS.n1306 1.5005
R4072 VSS.n1341 VSS.n1307 1.5005
R4073 VSS.n1441 VSS.n1311 1.5005
R4074 VSS.n1440 VSS.n1313 1.5005
R4075 VSS.n1439 VSS.n1315 1.5005
R4076 VSS.n1346 VSS.n1316 1.5005
R4077 VSS.n1435 VSS.n1320 1.5005
R4078 VSS.n1434 VSS.n1322 1.5005
R4079 VSS.n1433 VSS.n1324 1.5005
R4080 VSS.n1350 VSS.n1325 1.5005
R4081 VSS.n1429 VSS.n1329 1.5005
R4082 VSS.n1428 VSS.n1331 1.5005
R4083 VSS.n1427 VSS.n1333 1.5005
R4084 VSS.n1424 VSS.n1423 1.5005
R4085 VSS.n1422 VSS.n1421 1.5005
R4086 VSS.n3010 VSS.n2891 1.5005
R4087 VSS.n3012 VSS.n3011 1.5005
R4088 VSS.n3013 VSS.n2890 1.5005
R4089 VSS.n3015 VSS.n3014 1.5005
R4090 VSS.n3016 VSS.n2889 1.5005
R4091 VSS.n3018 VSS.n3017 1.5005
R4092 VSS.n3019 VSS.n2888 1.5005
R4093 VSS.n3021 VSS.n3020 1.5005
R4094 VSS.n3022 VSS.n2887 1.5005
R4095 VSS.n3024 VSS.n3023 1.5005
R4096 VSS.n3025 VSS.n2886 1.5005
R4097 VSS.n3027 VSS.n3026 1.5005
R4098 VSS.n3028 VSS.n2885 1.5005
R4099 VSS.n3030 VSS.n3029 1.5005
R4100 VSS.n3031 VSS.n2884 1.5005
R4101 VSS.n3033 VSS.n3032 1.5005
R4102 VSS.n3034 VSS.n2883 1.5005
R4103 VSS.n3036 VSS.n3035 1.5005
R4104 VSS.n3037 VSS.n2882 1.5005
R4105 VSS.n3039 VSS.n3038 1.5005
R4106 VSS.n1817 VSS.n897 1.45165
R4107 VSS.n1709 VSS.n936 1.45008
R4108 VSS.n1079 VSS.n1078 1.39283
R4109 VSS.n3232 VSS.n116 1.33629
R4110 VSS.n3251 VSS.n114 1.33629
R4111 VSS.n3251 VSS.n3250 1.33629
R4112 VSS.n3197 VSS.n3196 1.33629
R4113 VSS.n141 VSS.n102 1.33034
R4114 VSS.n1117 VSS.n1109 1.32992
R4115 VSS.n1117 VSS.n1108 1.32992
R4116 VSS.n1724 VSS.n1723 1.28295
R4117 VSS.n8 VSS.n0 1.2567
R4118 VSS.n901 VSS.n0 1.25289
R4119 VSS.n1817 VSS.n894 1.18996
R4120 VSS.n1835 VSS.n894 1.18996
R4121 VSS.n1835 VSS.n895 1.18996
R4122 VSS.n1831 VSS.n895 1.18996
R4123 VSS.n1831 VSS.n1821 1.18996
R4124 VSS.n1827 VSS.n1821 1.18996
R4125 VSS.n1827 VSS.n1824 1.18996
R4126 VSS.n1824 VSS.n1823 1.18996
R4127 VSS.n3425 VSS.n6 1.18996
R4128 VSS.n3420 VSS.n6 1.18996
R4129 VSS.n3420 VSS.n11 1.18996
R4130 VSS.n3416 VSS.n11 1.18996
R4131 VSS.n3416 VSS.n14 1.18996
R4132 VSS.n3412 VSS.n14 1.18996
R4133 VSS.n3412 VSS.n16 1.18996
R4134 VSS.n3408 VSS.n16 1.18996
R4135 VSS.n3408 VSS.n18 1.18996
R4136 VSS.n1553 VSS.n991 1.16769
R4137 VSS.n1334 VSS.n1332 1.16259
R4138 VSS.n3245 VSS.n117 1.16216
R4139 VSS.n187 VSS.n185 1.1255
R4140 VSS.n3112 VSS.n3111 1.1255
R4141 VSS.n3110 VSS.n186 1.1255
R4142 VSS.n3109 VSS.n3108 1.1255
R4143 VSS.n2834 VSS.n2828 1.1255
R4144 VSS.n2835 VSS.n2832 1.1255
R4145 VSS.n3100 VSS.n3099 1.1255
R4146 VSS.n3098 VSS.n2833 1.1255
R4147 VSS.n3097 VSS.n3096 1.1255
R4148 VSS.n2837 VSS.n2836 1.1255
R4149 VSS.n3090 VSS.n3089 1.1255
R4150 VSS.n3088 VSS.n2840 1.1255
R4151 VSS.n3087 VSS.n3086 1.1255
R4152 VSS.n2843 VSS.n2842 1.1255
R4153 VSS.n3080 VSS.n3079 1.1255
R4154 VSS.n3078 VSS.n2847 1.1255
R4155 VSS.n3077 VSS.n3076 1.1255
R4156 VSS.n2854 VSS.n2848 1.1255
R4157 VSS.n3070 VSS.n3069 1.1255
R4158 VSS.n3068 VSS.n2853 1.1255
R4159 VSS.n3067 VSS.n3066 1.1255
R4160 VSS.n2856 VSS.n2855 1.1255
R4161 VSS.n2870 VSS.n2858 1.1255
R4162 VSS.n2863 VSS.n2861 1.1255
R4163 VSS.n3056 VSS.n3055 1.1255
R4164 VSS.n3054 VSS.n2862 1.1255
R4165 VSS.n3053 VSS.n3052 1.1255
R4166 VSS.n2865 VSS.n2864 1.1255
R4167 VSS.n3046 VSS.n3045 1.1255
R4168 VSS.n3044 VSS.n2868 1.1255
R4169 VSS.n2922 VSS.n2869 1.1255
R4170 VSS.n2921 VSS.n2920 1.1255
R4171 VSS.n2917 VSS.n2916 1.1255
R4172 VSS.n2934 VSS.n2933 1.1255
R4173 VSS.n2935 VSS.n2915 1.1255
R4174 VSS.n2937 VSS.n2936 1.1255
R4175 VSS.n2938 VSS.n2872 1.1255
R4176 VSS.n2912 VSS.n2873 1.1255
R4177 VSS.n2946 VSS.n2945 1.1255
R4178 VSS.n2947 VSS.n2911 1.1255
R4179 VSS.n2950 VSS.n2949 1.1255
R4180 VSS.n2948 VSS.n2908 1.1255
R4181 VSS.n2956 VSS.n2874 1.1255
R4182 VSS.n2957 VSS.n2875 1.1255
R4183 VSS.n2963 VSS.n2962 1.1255
R4184 VSS.n2961 VSS.n2958 1.1255
R4185 VSS.n2960 VSS.n2905 1.1255
R4186 VSS.n2959 VSS.n2902 1.1255
R4187 VSS.n2974 VSS.n2903 1.1255
R4188 VSS.n2975 VSS.n2876 1.1255
R4189 VSS.n2976 VSS.n2877 1.1255
R4190 VSS.n2899 VSS.n2898 1.1255
R4191 VSS.n2984 VSS.n2983 1.1255
R4192 VSS.n2985 VSS.n2897 1.1255
R4193 VSS.n2987 VSS.n2986 1.1255
R4194 VSS.n2894 VSS.n2879 1.1255
R4195 VSS.n2994 VSS.n2880 1.1255
R4196 VSS.n2997 VSS.n2995 1.1255
R4197 VSS.n3000 VSS.n2999 1.1255
R4198 VSS.n2998 VSS.n2996 1.1255
R4199 VSS.n2881 VSS.n2878 1.1255
R4200 VSS.n2827 VSS.n2826 1.1255
R4201 VSS.n185 VSS.n183 1.1255
R4202 VSS.n3113 VSS.n3112 1.1255
R4203 VSS.n186 VSS.n184 1.1255
R4204 VSS.n3108 VSS.n3107 1.1255
R4205 VSS.n3105 VSS.n2828 1.1255
R4206 VSS.n2832 VSS.n2829 1.1255
R4207 VSS.n3101 VSS.n3100 1.1255
R4208 VSS.n2833 VSS.n2831 1.1255
R4209 VSS.n3096 VSS.n3095 1.1255
R4210 VSS.n2838 VSS.n2837 1.1255
R4211 VSS.n3091 VSS.n3090 1.1255
R4212 VSS.n2840 VSS.n2839 1.1255
R4213 VSS.n3086 VSS.n3085 1.1255
R4214 VSS.n2844 VSS.n2843 1.1255
R4215 VSS.n3081 VSS.n3080 1.1255
R4216 VSS.n2847 VSS.n2846 1.1255
R4217 VSS.n3076 VSS.n3075 1.1255
R4218 VSS.n2849 VSS.n2848 1.1255
R4219 VSS.n3071 VSS.n3070 1.1255
R4220 VSS.n2853 VSS.n2852 1.1255
R4221 VSS.n3066 VSS.n3065 1.1255
R4222 VSS.n3062 VSS.n2856 1.1255
R4223 VSS.n3061 VSS.n2858 1.1255
R4224 VSS.n2861 VSS.n2857 1.1255
R4225 VSS.n3057 VSS.n3056 1.1255
R4226 VSS.n2862 VSS.n2860 1.1255
R4227 VSS.n3052 VSS.n3051 1.1255
R4228 VSS.n2866 VSS.n2865 1.1255
R4229 VSS.n3047 VSS.n3046 1.1255
R4230 VSS.n2868 VSS.n2867 1.1255
R4231 VSS.n2923 VSS.n2922 1.1255
R4232 VSS.n2921 VSS.n2918 1.1255
R4233 VSS.n2927 VSS.n2917 1.1255
R4234 VSS.n2933 VSS.n2932 1.1255
R4235 VSS.n2928 VSS.n2915 1.1255
R4236 VSS.n2937 VSS.n2914 1.1255
R4237 VSS.n2939 VSS.n2938 1.1255
R4238 VSS.n2913 VSS.n2912 1.1255
R4239 VSS.n2945 VSS.n2944 1.1255
R4240 VSS.n2911 VSS.n2910 1.1255
R4241 VSS.n2951 VSS.n2950 1.1255
R4242 VSS.n2909 VSS.n2908 1.1255
R4243 VSS.n2956 VSS.n2955 1.1255
R4244 VSS.n2957 VSS.n2907 1.1255
R4245 VSS.n2964 VSS.n2963 1.1255
R4246 VSS.n2958 VSS.n2904 1.1255
R4247 VSS.n2968 VSS.n2905 1.1255
R4248 VSS.n2969 VSS.n2902 1.1255
R4249 VSS.n2974 VSS.n2973 1.1255
R4250 VSS.n2975 VSS.n2901 1.1255
R4251 VSS.n2977 VSS.n2976 1.1255
R4252 VSS.n2900 VSS.n2899 1.1255
R4253 VSS.n2983 VSS.n2982 1.1255
R4254 VSS.n2897 VSS.n2896 1.1255
R4255 VSS.n2988 VSS.n2987 1.1255
R4256 VSS.n2895 VSS.n2894 1.1255
R4257 VSS.n2994 VSS.n2993 1.1255
R4258 VSS.n2995 VSS.n2893 1.1255
R4259 VSS.n3001 VSS.n3000 1.1255
R4260 VSS.n2996 VSS.n2892 1.1255
R4261 VSS.n3005 VSS.n2881 1.1255
R4262 VSS.n2826 VSS.n2825 1.1255
R4263 VSS.n3005 VSS.n3004 1.1255
R4264 VSS.n3003 VSS.n2892 1.1255
R4265 VSS.n3002 VSS.n3001 1.1255
R4266 VSS.n2991 VSS.n2893 1.1255
R4267 VSS.n2993 VSS.n2992 1.1255
R4268 VSS.n2990 VSS.n2895 1.1255
R4269 VSS.n2989 VSS.n2988 1.1255
R4270 VSS.n2980 VSS.n2896 1.1255
R4271 VSS.n2982 VSS.n2981 1.1255
R4272 VSS.n2979 VSS.n2900 1.1255
R4273 VSS.n2978 VSS.n2977 1.1255
R4274 VSS.n2971 VSS.n2901 1.1255
R4275 VSS.n2973 VSS.n2972 1.1255
R4276 VSS.n2970 VSS.n2969 1.1255
R4277 VSS.n2968 VSS.n2967 1.1255
R4278 VSS.n2966 VSS.n2904 1.1255
R4279 VSS.n2965 VSS.n2964 1.1255
R4280 VSS.n2907 VSS.n2906 1.1255
R4281 VSS.n2955 VSS.n2954 1.1255
R4282 VSS.n2953 VSS.n2909 1.1255
R4283 VSS.n2952 VSS.n2951 1.1255
R4284 VSS.n2942 VSS.n2910 1.1255
R4285 VSS.n2944 VSS.n2943 1.1255
R4286 VSS.n2941 VSS.n2913 1.1255
R4287 VSS.n2940 VSS.n2939 1.1255
R4288 VSS.n2929 VSS.n2914 1.1255
R4289 VSS.n2930 VSS.n2928 1.1255
R4290 VSS.n2932 VSS.n2931 1.1255
R4291 VSS.n2927 VSS.n2926 1.1255
R4292 VSS.n2925 VSS.n2918 1.1255
R4293 VSS.n2924 VSS.n2923 1.1255
R4294 VSS.n2919 VSS.n2867 1.1255
R4295 VSS.n3048 VSS.n3047 1.1255
R4296 VSS.n3049 VSS.n2866 1.1255
R4297 VSS.n3051 VSS.n3050 1.1255
R4298 VSS.n2860 VSS.n2859 1.1255
R4299 VSS.n3058 VSS.n3057 1.1255
R4300 VSS.n3059 VSS.n2857 1.1255
R4301 VSS.n3061 VSS.n3060 1.1255
R4302 VSS.n3063 VSS.n3062 1.1255
R4303 VSS.n3065 VSS.n3064 1.1255
R4304 VSS.n2852 VSS.n2851 1.1255
R4305 VSS.n3072 VSS.n3071 1.1255
R4306 VSS.n3073 VSS.n2849 1.1255
R4307 VSS.n3075 VSS.n3074 1.1255
R4308 VSS.n2850 VSS.n2846 1.1255
R4309 VSS.n3082 VSS.n3081 1.1255
R4310 VSS.n3083 VSS.n2844 1.1255
R4311 VSS.n3085 VSS.n3084 1.1255
R4312 VSS.n2845 VSS.n2839 1.1255
R4313 VSS.n3092 VSS.n3091 1.1255
R4314 VSS.n3093 VSS.n2838 1.1255
R4315 VSS.n3095 VSS.n3094 1.1255
R4316 VSS.n2831 VSS.n2830 1.1255
R4317 VSS.n3102 VSS.n3101 1.1255
R4318 VSS.n3103 VSS.n2829 1.1255
R4319 VSS.n3105 VSS.n3104 1.1255
R4320 VSS.n3107 VSS.n3106 1.1255
R4321 VSS.n184 VSS.n182 1.1255
R4322 VSS.n3114 VSS.n3113 1.1255
R4323 VSS.n183 VSS.n181 1.1255
R4324 VSS.n2825 VSS.n2824 1.1255
R4325 VSS.n991 VSS.n907 1.0535
R4326 VSS.n3423 VSS.n9 1.05237
R4327 VSS.n1078 VSS.n906 0.977
R4328 VSS.n3228 VSS.n120 0.94832
R4329 VSS.n1923 VSS.n1922 0.939203
R4330 VSS.n1923 VSS.n812 0.939203
R4331 VSS.n2026 VSS.n785 0.939203
R4332 VSS.n2029 VSS.n785 0.939203
R4333 VSS.n2200 VSS.n2199 0.939203
R4334 VSS.n2200 VSS.n633 0.939203
R4335 VSS.n2303 VSS.n606 0.939203
R4336 VSS.n2306 VSS.n606 0.939203
R4337 VSS.n2527 VSS.n456 0.939203
R4338 VSS.n2527 VSS.n454 0.939203
R4339 VSS.n2338 VSS.n543 0.939203
R4340 VSS.n2338 VSS.n542 0.939203
R4341 VSS.n2489 VSS.n2488 0.939203
R4342 VSS.n2489 VSS.n476 0.939203
R4343 VSS.n2749 VSS.n259 0.939203
R4344 VSS.n259 VSS.n258 0.939203
R4345 VSS.n1886 VSS.n1885 0.939203
R4346 VSS.n1886 VSS.n831 0.939203
R4347 VSS.n2061 VSS.n722 0.939203
R4348 VSS.n2061 VSS.n721 0.939203
R4349 VSS.n2163 VSS.n652 0.939203
R4350 VSS.n2163 VSS.n2162 0.939203
R4351 VSS.n2338 VSS.n541 0.939203
R4352 VSS.n2338 VSS.n540 0.939203
R4353 VSS.n2490 VSS.n2489 0.939203
R4354 VSS.n2489 VSS.n475 0.939203
R4355 VSS.n2163 VSS.n651 0.939203
R4356 VSS.n2163 VSS.n650 0.939203
R4357 VSS.n685 VSS.n684 0.939203
R4358 VSS.n684 VSS.n657 0.939203
R4359 VSS.n684 VSS.n658 0.939203
R4360 VSS.n684 VSS.n659 0.939203
R4361 VSS.n577 VSS.n576 0.939203
R4362 VSS.n576 VSS.n549 0.939203
R4363 VSS.n576 VSS.n550 0.939203
R4364 VSS.n576 VSS.n551 0.939203
R4365 VSS.n507 VSS.n193 0.939203
R4366 VSS.n501 VSS.n193 0.939203
R4367 VSS.n499 VSS.n193 0.939203
R4368 VSS.n493 VSS.n193 0.939203
R4369 VSS.n2756 VSS.n251 0.939203
R4370 VSS.n255 VSS.n251 0.939203
R4371 VSS.n2763 VSS.n251 0.939203
R4372 VSS.n2766 VSS.n251 0.939203
R4373 VSS.n2579 VSS.n422 0.939203
R4374 VSS.n426 VSS.n422 0.939203
R4375 VSS.n2406 VSS.n259 0.939203
R4376 VSS.n2404 VSS.n259 0.939203
R4377 VSS.n2061 VSS.n720 0.939203
R4378 VSS.n2061 VSS.n719 0.939203
R4379 VSS.n756 VSS.n755 0.939203
R4380 VSS.n755 VSS.n728 0.939203
R4381 VSS.n755 VSS.n729 0.939203
R4382 VSS.n755 VSS.n730 0.939203
R4383 VSS.n348 VSS.n286 0.939203
R4384 VSS.n342 VSS.n286 0.939203
R4385 VSS.n340 VSS.n286 0.939203
R4386 VSS.n334 VSS.n286 0.939203
R4387 VSS.n329 VSS.n328 0.939203
R4388 VSS.n2650 VSS.n2649 0.939203
R4389 VSS.n2650 VSS.n2625 0.939203
R4390 VSS.n2650 VSS.n2624 0.939203
R4391 VSS.n2650 VSS.n2623 0.939203
R4392 VSS.n355 VSS.n286 0.939203
R4393 VSS.n354 VSS.n286 0.939203
R4394 VSS.n362 VSS.n286 0.939203
R4395 VSS.n365 VSS.n286 0.939203
R4396 VSS.n140 VSS.n130 0.939203
R4397 VSS.n3212 VSS.n130 0.939203
R4398 VSS.n3215 VSS.n130 0.939203
R4399 VSS.n2732 VSS.n268 0.939203
R4400 VSS.n2735 VSS.n268 0.939203
R4401 VSS.n1886 VSS.n830 0.939203
R4402 VSS.n1886 VSS.n829 0.939203
R4403 VSS.n1867 VSS.n1866 0.939203
R4404 VSS.n1866 VSS.n1838 0.939203
R4405 VSS.n1866 VSS.n1839 0.939203
R4406 VSS.n1866 VSS.n1840 0.939203
R4407 VSS.n1848 VSS.n1847 0.939203
R4408 VSS.n1847 VSS.n1846 0.939203
R4409 VSS.n737 VSS.n40 0.939203
R4410 VSS.n735 VSS.n40 0.939203
R4411 VSS.n666 VSS.n62 0.939203
R4412 VSS.n664 VSS.n62 0.939203
R4413 VSS.n558 VSS.n84 0.939203
R4414 VSS.n556 VSS.n84 0.939203
R4415 VSS.n2821 VSS.n190 0.939203
R4416 VSS.n2821 VSS.n189 0.939203
R4417 VSS.n2780 VSS.n2772 0.939203
R4418 VSS.n2780 VSS.n242 0.939203
R4419 VSS.n3119 VSS.n98 0.939203
R4420 VSS.n3126 VSS.n98 0.939203
R4421 VSS.n3132 VSS.n100 0.939203
R4422 VSS.n3135 VSS.n100 0.939203
R4423 VSS.n3141 VSS.n100 0.939203
R4424 VSS.n3144 VSS.n100 0.939203
R4425 VSS.n3150 VSS.n100 0.939203
R4426 VSS.n3152 VSS.n100 0.939203
R4427 VSS.n3158 VSS.n100 0.939203
R4428 VSS.n3160 VSS.n100 0.939203
R4429 VSS.n3166 VSS.n100 0.939203
R4430 VSS.n3168 VSS.n100 0.939203
R4431 VSS.n3174 VSS.n100 0.939203
R4432 VSS.n3176 VSS.n100 0.939203
R4433 VSS.n3182 VSS.n100 0.939203
R4434 VSS.n1616 VSS.n933 0.93088
R4435 VSS.n1231 VSS.n1229 0.9185
R4436 VSS.n411 VSS.n410 0.915775
R4437 VSS.n3186 VSS.n107 0.907605
R4438 VSS.n1823 VSS.n3 0.904493
R4439 VSS.n3008 VSS.n3007 0.9005
R4440 VSS.n3228 VSS.n3227 0.871619
R4441 VSS.n3190 VSS.n115 0.867167
R4442 VSS.n3193 VSS.n3192 0.867167
R4443 VSS.n3192 VSS.n110 0.867167
R4444 VSS.n1420 VSS.t43 0.833115
R4445 VSS.n2633 VSS.t137 0.8195
R4446 VSS.n2633 VSS.t246 0.8195
R4447 VSS.n2634 VSS.t161 0.8195
R4448 VSS.n2634 VSS.t131 0.8195
R4449 VSS.n1725 VSS.n1724 0.807125
R4450 VSS.n1186 VSS.n1072 0.779896
R4451 VSS.t209 VSS.n2827 0.758022
R4452 VSS.n3196 VSS.n3195 0.73471
R4453 VSS.n1198 VSS.n1197 0.705167
R4454 VSS.n1198 VSS.n1087 0.705167
R4455 VSS.n1198 VSS.n1088 0.705167
R4456 VSS.n1198 VSS.n1089 0.705167
R4457 VSS.n1198 VSS.n1090 0.705167
R4458 VSS.n1198 VSS.n1091 0.705167
R4459 VSS.n1198 VSS.n1092 0.705167
R4460 VSS.n1198 VSS.n1093 0.705167
R4461 VSS.n1032 VSS.n1017 0.705167
R4462 VSS.n1038 VSS.n1017 0.705167
R4463 VSS.n1030 VSS.n1017 0.705167
R4464 VSS.n1045 VSS.n1017 0.705167
R4465 VSS.n1027 VSS.n1017 0.705167
R4466 VSS.n1052 VSS.n1017 0.705167
R4467 VSS.n1024 VSS.n1017 0.705167
R4468 VSS.n1059 VSS.n1017 0.705167
R4469 VSS.n1550 VSS.n995 0.698475
R4470 VSS.n1550 VSS.n996 0.698475
R4471 VSS.n1550 VSS.n997 0.698475
R4472 VSS.n1550 VSS.n998 0.698475
R4473 VSS.n1550 VSS.n999 0.698475
R4474 VSS.n1550 VSS.n1000 0.698475
R4475 VSS.n1550 VSS.n1001 0.698475
R4476 VSS.n1705 VSS.n1704 0.690672
R4477 VSS.n1656 VSS.n1633 0.660831
R4478 VSS.n1945 VSS.n1944 0.660831
R4479 VSS.n1979 VSS.n1978 0.660831
R4480 VSS.n2222 VSS.n2221 0.660831
R4481 VSS.n2256 VSS.n2255 0.660831
R4482 VSS.n2549 VSS.n440 0.660831
R4483 VSS.n3041 VSS.n2881 0.64962
R4484 VSS.n21 VSS.n18 0.642811
R4485 VSS.n1709 VSS.n1708 0.608375
R4486 VSS.n1708 VSS.n1707 0.608
R4487 VSS.n1450 VSS.n9 0.58325
R4488 VSS.n3187 VSS.n3185 0.567737
R4489 VSS.n3208 VSS.n139 0.553526
R4490 VSS.n1518 VSS.n1005 0.545237
R4491 VSS.n1550 VSS.n994 0.538771
R4492 VSS.n1726 VSS.n925 0.532146
R4493 VSS.n1519 VSS.n1518 0.513263
R4494 VSS.n1471 VSS.n1470 0.50099
R4495 VSS.n1465 VSS.n1286 0.5005
R4496 VSS.n1363 VSS.n1255 0.5005
R4497 VSS.n1375 VSS.n1257 0.5005
R4498 VSS.n1362 VSS.n1254 0.5005
R4499 VSS.n1376 VSS.n1258 0.5005
R4500 VSS.n1361 VSS.n1253 0.5005
R4501 VSS.n1377 VSS.n1259 0.5005
R4502 VSS.n1360 VSS.n1252 0.5005
R4503 VSS.n1378 VSS.n1260 0.5005
R4504 VSS.n1359 VSS.n1251 0.5005
R4505 VSS.n1379 VSS.n1261 0.5005
R4506 VSS.n1358 VSS.n1250 0.5005
R4507 VSS.n1380 VSS.n1262 0.5005
R4508 VSS.n1357 VSS.n1249 0.5005
R4509 VSS.n1381 VSS.n1263 0.5005
R4510 VSS.n1356 VSS.n1248 0.5005
R4511 VSS.n1417 VSS.n1264 0.5005
R4512 VSS.n1382 VSS.n1247 0.5005
R4513 VSS.n1467 VSS.n1268 0.5005
R4514 VSS.n1454 VSS.n1291 0.5005
R4515 VSS.n1374 VSS.n1295 0.5005
R4516 VSS.n1372 VSS.n1371 0.5005
R4517 VSS.n1706 VSS.n1705 0.4835
R4518 VSS.n1034 VSS.n1015 0.476553
R4519 VSS.n1063 VSS.n1062 0.471816
R4520 VSS.n1469 VSS.n1245 0.460063
R4521 VSS.n3197 VSS.n3193 0.458789
R4522 VSS.n3193 VSS.n114 0.458789
R4523 VSS.n3009 VSS.n105 0.451478
R4524 VSS.n1241 VSS.n1240 0.43349
R4525 VSS.n1086 VSS.n1073 0.419711
R4526 VSS.n3250 VSS.n115 0.413789
R4527 VSS.n1153 VSS.n1083 0.4082
R4528 VSS.n1078 VSS.n2 0.4005
R4529 VSS.n898 VSS.n2 0.4005
R4530 VSS.n3244 VSS.n3243 0.394162
R4531 VSS.n1472 VSS.n1243 0.39128
R4532 VSS.n1199 VSS.n1086 0.3866
R4533 VSS.n1203 VSS.n1082 0.3668
R4534 VSS.n1547 VSS.n1546 0.365237
R4535 VSS.n1546 VSS.n1543 0.365237
R4536 VSS.n1543 VSS.n1542 0.365237
R4537 VSS.n1542 VSS.n1539 0.365237
R4538 VSS.n1539 VSS.n1538 0.365237
R4539 VSS.n1538 VSS.n1535 0.365237
R4540 VSS.n1535 VSS.n1534 0.365237
R4541 VSS.n1534 VSS.n1531 0.365237
R4542 VSS.n1531 VSS.n1530 0.365237
R4543 VSS.n1530 VSS.n1527 0.365237
R4544 VSS.n1527 VSS.n1526 0.365237
R4545 VSS.n1526 VSS.n1523 0.365237
R4546 VSS.n1523 VSS.n1522 0.365237
R4547 VSS.n1522 VSS.n1519 0.365237
R4548 VSS.n1125 VSS.n1124 0.3605
R4549 VSS.n1127 VSS.n1125 0.3605
R4550 VSS.n1128 VSS.n1127 0.3605
R4551 VSS.n1131 VSS.n1128 0.3605
R4552 VSS.n1132 VSS.n1131 0.3605
R4553 VSS.n1135 VSS.n1132 0.3605
R4554 VSS.n1136 VSS.n1135 0.3605
R4555 VSS.n1139 VSS.n1136 0.3605
R4556 VSS.n1140 VSS.n1139 0.3605
R4557 VSS.n1143 VSS.n1140 0.3605
R4558 VSS.n1144 VSS.n1143 0.3605
R4559 VSS.n1147 VSS.n1144 0.3605
R4560 VSS.n1148 VSS.n1147 0.3605
R4561 VSS.n1151 VSS.n1148 0.3605
R4562 VSS.n1154 VSS.n1151 0.3605
R4563 VSS.n1085 VSS.n1074 0.3605
R4564 VSS.n1200 VSS.n1085 0.3605
R4565 VSS.n1200 VSS.n1199 0.3605
R4566 VSS.n1062 VSS.n1021 0.3605
R4567 VSS.n1057 VSS.n1021 0.3605
R4568 VSS.n1057 VSS.n1056 0.3605
R4569 VSS.n1056 VSS.n1055 0.3605
R4570 VSS.n1055 VSS.n1023 0.3605
R4571 VSS.n1050 VSS.n1023 0.3605
R4572 VSS.n1050 VSS.n1049 0.3605
R4573 VSS.n1049 VSS.n1048 0.3605
R4574 VSS.n1048 VSS.n1026 0.3605
R4575 VSS.n1043 VSS.n1026 0.3605
R4576 VSS.n1043 VSS.n1042 0.3605
R4577 VSS.n1042 VSS.n1041 0.3605
R4578 VSS.n1041 VSS.n1029 0.3605
R4579 VSS.n1036 VSS.n1029 0.3605
R4580 VSS.n1036 VSS.n1035 0.3605
R4581 VSS.n1035 VSS.n1034 0.3605
R4582 VSS.n1203 VSS.n1202 0.3578
R4583 VSS.n1202 VSS.n1083 0.3461
R4584 VSS.n1208 VSS.n1207 0.3317
R4585 VSS.n1207 VSS.n965 0.3317
R4586 VSS.n1559 VSS.n1558 0.3317
R4587 VSS.n1194 VSS.n1193 0.313132
R4588 VSS.n1193 VSS.n1192 0.313132
R4589 VSS.n1192 VSS.n1098 0.313132
R4590 VSS.n1158 VSS.n1123 0.313132
R4591 VSS.n1159 VSS.n1158 0.313132
R4592 VSS.n1160 VSS.n1159 0.313132
R4593 VSS.n1161 VSS.n1160 0.313132
R4594 VSS.n1162 VSS.n1161 0.313132
R4595 VSS.n1163 VSS.n1162 0.313132
R4596 VSS.n1164 VSS.n1163 0.313132
R4597 VSS.n1166 VSS.n1164 0.313132
R4598 VSS.n1167 VSS.n1166 0.313132
R4599 VSS.n1168 VSS.n1167 0.313132
R4600 VSS.n1497 VSS.n1496 0.313132
R4601 VSS.n1498 VSS.n1497 0.313132
R4602 VSS.n1498 VSS.n1011 0.313132
R4603 VSS.n1504 VSS.n1011 0.313132
R4604 VSS.n1505 VSS.n1504 0.313132
R4605 VSS.n1506 VSS.n1505 0.313132
R4606 VSS.n1506 VSS.n1007 0.313132
R4607 VSS.n1513 VSS.n1007 0.313132
R4608 VSS.n1514 VSS.n1513 0.313132
R4609 VSS.n1515 VSS.n1514 0.313132
R4610 VSS.n1175 VSS.n1174 0.313132
R4611 VSS.n1174 VSS.n1173 0.313132
R4612 VSS.n1173 VSS.n1119 0.313132
R4613 VSS.n1492 VSS.n1491 0.313132
R4614 VSS.n1491 VSS.n1490 0.313132
R4615 VSS.n1490 VSS.n1064 0.313132
R4616 VSS.n1484 VSS.n1064 0.313132
R4617 VSS.n1484 VSS.n1483 0.313132
R4618 VSS.n1483 VSS.n1482 0.313132
R4619 VSS.n1482 VSS.n1068 0.313132
R4620 VSS.n1476 VSS.n1068 0.313132
R4621 VSS.n1476 VSS.n1475 0.313132
R4622 VSS.n1475 VSS.n1474 0.313132
R4623 VSS.n1118 VSS.n1098 0.311947
R4624 VSS.n1548 VSS.n1547 0.311947
R4625 VSS.n1152 VSS.n1077 0.310763
R4626 VSS.n1079 VSS.n1005 0.310763
R4627 VSS.n1080 VSS.n1079 0.3015
R4628 VSS.n1124 VSS.n1086 0.294184
R4629 VSS.n1710 VSS.n1709 0.289389
R4630 VSS.n1553 VSS.n1552 0.289389
R4631 VSS.n1552 VSS.n1551 0.289389
R4632 VSS.n1711 VSS.n1710 0.289181
R4633 VSS.n1692 VSS.n1691 0.286527
R4634 VSS.n1691 VSS.n1690 0.286527
R4635 VSS.n1241 VSS.n1074 0.2849
R4636 VSS.n1242 VSS.n1241 0.27473
R4637 VSS.n1240 VSS.n1075 0.2741
R4638 VSS.n1239 VSS.n1076 0.2705
R4639 VSS.n1175 VSS.n1118 0.2705
R4640 VSS.n1725 VSS.n926 0.269375
R4641 VSS.n3265 VSS.n3264 0.265655
R4642 VSS.n1245 VSS.n8 0.254021
R4643 VSS.n1812 VSS.n1811 0.254021
R4644 VSS.n1811 VSS.n1810 0.254021
R4645 VSS.n1810 VSS.n1808 0.254021
R4646 VSS.n1808 VSS.n902 0.254021
R4647 VSS.n1803 VSS.n902 0.254021
R4648 VSS.n1803 VSS.n1802 0.254021
R4649 VSS.n1802 VSS.n1801 0.254021
R4650 VSS.n1795 VSS.n908 0.254021
R4651 VSS.n1790 VSS.n908 0.254021
R4652 VSS.n1790 VSS.n1789 0.254021
R4653 VSS.n1789 VSS.n1788 0.254021
R4654 VSS.n1788 VSS.n910 0.254021
R4655 VSS.n921 VSS.n910 0.254021
R4656 VSS.n923 VSS.n921 0.254021
R4657 VSS.n1730 VSS.n1728 0.254021
R4658 VSS.n1728 VSS.n924 0.254021
R4659 VSS.n1588 VSS.n924 0.254021
R4660 VSS.n1592 VSS.n1588 0.254021
R4661 VSS.n1593 VSS.n1592 0.254021
R4662 VSS.n1594 VSS.n1593 0.254021
R4663 VSS.n1594 VSS.n1584 0.254021
R4664 VSS.n1601 VSS.n1584 0.254021
R4665 VSS.n1602 VSS.n1601 0.254021
R4666 VSS.n1603 VSS.n1602 0.254021
R4667 VSS.n1607 VSS.n1606 0.254021
R4668 VSS.n1608 VSS.n1607 0.254021
R4669 VSS.n1608 VSS.n1579 0.254021
R4670 VSS.n1614 VSS.n1579 0.254021
R4671 VSS.n1615 VSS.n1614 0.254021
R4672 VSS.n1623 VSS.n1615 0.254021
R4673 VSS.n1623 VSS.n1622 0.254021
R4674 VSS.n1622 VSS.n1621 0.254021
R4675 VSS.n1621 VSS.n1618 0.254021
R4676 VSS.n1618 VSS.n1617 0.254021
R4677 VSS.n3252 VSS.n3251 0.248119
R4678 VSS.t201 VSS.n3252 0.248119
R4679 VSS.n1237 VSS.n1236 0.248119
R4680 VSS.n1236 VSS.n1235 0.248119
R4681 VSS.n1707 VSS.n939 0.243993
R4682 VSS.n1705 VSS.n1697 0.243993
R4683 VSS.n1233 VSS.n936 0.2408
R4684 VSS.n3426 VSS.n3 0.238393
R4685 VSS.n1843 VSS.n19 0.237342
R4686 VSS.n1850 VSS.n1843 0.237342
R4687 VSS.n1851 VSS.n1850 0.237342
R4688 VSS.n1864 VSS.n1851 0.237342
R4689 VSS.n1864 VSS.n1863 0.237342
R4690 VSS.n1863 VSS.n1862 0.237342
R4691 VSS.n1862 VSS.n1859 0.237342
R4692 VSS.n1859 VSS.n1858 0.237342
R4693 VSS.n1858 VSS.n1855 0.237342
R4694 VSS.n1855 VSS.n1854 0.237342
R4695 VSS.n1854 VSS.n1852 0.237342
R4696 VSS.n1852 VSS.n887 0.237342
R4697 VSS.n1870 VSS.n887 0.237342
R4698 VSS.n1871 VSS.n1870 0.237342
R4699 VSS.n1874 VSS.n1871 0.237342
R4700 VSS.n1875 VSS.n1874 0.237342
R4701 VSS.n316 VSS.n153 0.237342
R4702 VSS.n317 VSS.n316 0.237342
R4703 VSS.n317 VSS.n310 0.237342
R4704 VSS.n323 VSS.n310 0.237342
R4705 VSS.n324 VSS.n323 0.237342
R4706 VSS.n326 VSS.n324 0.237342
R4707 VSS.n326 VSS.n325 0.237342
R4708 VSS.n325 VSS.n307 0.237342
R4709 VSS.n336 VSS.n307 0.237342
R4710 VSS.n337 VSS.n336 0.237342
R4711 VSS.n338 VSS.n337 0.237342
R4712 VSS.n338 VSS.n305 0.237342
R4713 VSS.n344 VSS.n305 0.237342
R4714 VSS.n345 VSS.n344 0.237342
R4715 VSS.n346 VSS.n345 0.237342
R4716 VSS.n346 VSS.n302 0.237342
R4717 VSS.n367 VSS.n303 0.237342
R4718 VSS.n351 VSS.n303 0.237342
R4719 VSS.n360 VSS.n351 0.237342
R4720 VSS.n360 VSS.n359 0.237342
R4721 VSS.n359 VSS.n358 0.237342
R4722 VSS.n358 VSS.n353 0.237342
R4723 VSS.n353 VSS.n290 0.237342
R4724 VSS.n2705 VSS.n290 0.237342
R4725 VSS.n2705 VSS.n2704 0.237342
R4726 VSS.n2704 VSS.n2703 0.237342
R4727 VSS.n2703 VSS.n291 0.237342
R4728 VSS.n2628 VSS.n291 0.237342
R4729 VSS.n2628 VSS.n2627 0.237342
R4730 VSS.n2640 VSS.n2637 0.237342
R4731 VSS.n2641 VSS.n2640 0.237342
R4732 VSS.n2644 VSS.n2641 0.237342
R4733 VSS.n2645 VSS.n2644 0.237342
R4734 VSS.n2646 VSS.n2645 0.237342
R4735 VSS.n2646 VSS.n400 0.237342
R4736 VSS.n248 VSS.n246 0.237342
R4737 VSS.n249 VSS.n248 0.237342
R4738 VSS.n2770 VSS.n249 0.237342
R4739 VSS.n2770 VSS.n2769 0.237342
R4740 VSS.n2769 VSS.n2768 0.237342
R4741 VSS.n2768 VSS.n250 0.237342
R4742 VSS.n252 VSS.n250 0.237342
R4743 VSS.n2761 VSS.n252 0.237342
R4744 VSS.n2761 VSS.n2760 0.237342
R4745 VSS.n2760 VSS.n2759 0.237342
R4746 VSS.n2759 VSS.n254 0.237342
R4747 VSS.n2754 VSS.n254 0.237342
R4748 VSS.n2754 VSS.n2753 0.237342
R4749 VSS.n2753 VSS.n2752 0.237342
R4750 VSS.n2752 VSS.n257 0.237342
R4751 VSS.n2747 VSS.n257 0.237342
R4752 VSS.n486 VSS.n485 0.237342
R4753 VSS.n489 VSS.n486 0.237342
R4754 VSS.n490 VSS.n489 0.237342
R4755 VSS.n490 VSS.n483 0.237342
R4756 VSS.n495 VSS.n483 0.237342
R4757 VSS.n496 VSS.n495 0.237342
R4758 VSS.n497 VSS.n496 0.237342
R4759 VSS.n497 VSS.n481 0.237342
R4760 VSS.n503 VSS.n481 0.237342
R4761 VSS.n504 VSS.n503 0.237342
R4762 VSS.n505 VSS.n504 0.237342
R4763 VSS.n505 VSS.n479 0.237342
R4764 VSS.n510 VSS.n479 0.237342
R4765 VSS.n512 VSS.n510 0.237342
R4766 VSS.n513 VSS.n512 0.237342
R4767 VSS.n2486 VSS.n513 0.237342
R4768 VSS.n554 VSS.n86 0.237342
R4769 VSS.n560 VSS.n554 0.237342
R4770 VSS.n561 VSS.n560 0.237342
R4771 VSS.n574 VSS.n561 0.237342
R4772 VSS.n574 VSS.n573 0.237342
R4773 VSS.n573 VSS.n572 0.237342
R4774 VSS.n572 VSS.n569 0.237342
R4775 VSS.n569 VSS.n568 0.237342
R4776 VSS.n568 VSS.n565 0.237342
R4777 VSS.n565 VSS.n564 0.237342
R4778 VSS.n564 VSS.n562 0.237342
R4779 VSS.n562 VSS.n547 0.237342
R4780 VSS.n580 VSS.n547 0.237342
R4781 VSS.n581 VSS.n580 0.237342
R4782 VSS.n584 VSS.n581 0.237342
R4783 VSS.n585 VSS.n584 0.237342
R4784 VSS.n1881 VSS.n1879 0.237342
R4785 VSS.n1882 VSS.n1881 0.237342
R4786 VSS.n1883 VSS.n1882 0.237342
R4787 VSS.n1883 VSS.n826 0.237342
R4788 VSS.n1891 VSS.n826 0.237342
R4789 VSS.n1892 VSS.n1891 0.237342
R4790 VSS.n1893 VSS.n1892 0.237342
R4791 VSS.n1893 VSS.n822 0.237342
R4792 VSS.n1899 VSS.n822 0.237342
R4793 VSS.n1900 VSS.n1899 0.237342
R4794 VSS.n1901 VSS.n1900 0.237342
R4795 VSS.n1901 VSS.n818 0.237342
R4796 VSS.n1907 VSS.n818 0.237342
R4797 VSS.n1908 VSS.n1907 0.237342
R4798 VSS.n1910 VSS.n1908 0.237342
R4799 VSS.n1910 VSS.n1909 0.237342
R4800 VSS.n1909 VSS.n814 0.237342
R4801 VSS.n1917 VSS.n814 0.237342
R4802 VSS.n1918 VSS.n1917 0.237342
R4803 VSS.n1919 VSS.n1918 0.237342
R4804 VSS.n1919 VSS.n808 0.237342
R4805 VSS.n767 VSS.n766 0.237342
R4806 VSS.n770 VSS.n767 0.237342
R4807 VSS.n771 VSS.n770 0.237342
R4808 VSS.n2057 VSS.n771 0.237342
R4809 VSS.n2057 VSS.n2056 0.237342
R4810 VSS.n2056 VSS.n2055 0.237342
R4811 VSS.n2055 VSS.n772 0.237342
R4812 VSS.n2049 VSS.n772 0.237342
R4813 VSS.n2049 VSS.n2048 0.237342
R4814 VSS.n2048 VSS.n2047 0.237342
R4815 VSS.n2047 VSS.n776 0.237342
R4816 VSS.n2041 VSS.n776 0.237342
R4817 VSS.n2041 VSS.n2040 0.237342
R4818 VSS.n2040 VSS.n2039 0.237342
R4819 VSS.n2039 VSS.n780 0.237342
R4820 VSS.n2033 VSS.n780 0.237342
R4821 VSS.n2033 VSS.n2032 0.237342
R4822 VSS.n2032 VSS.n2031 0.237342
R4823 VSS.n2031 VSS.n784 0.237342
R4824 VSS.n786 VSS.n784 0.237342
R4825 VSS.n2024 VSS.n786 0.237342
R4826 VSS.n2160 VSS.n2156 0.237342
R4827 VSS.n2160 VSS.n2159 0.237342
R4828 VSS.n2159 VSS.n2158 0.237342
R4829 VSS.n2158 VSS.n647 0.237342
R4830 VSS.n2168 VSS.n647 0.237342
R4831 VSS.n2169 VSS.n2168 0.237342
R4832 VSS.n2170 VSS.n2169 0.237342
R4833 VSS.n2170 VSS.n643 0.237342
R4834 VSS.n2176 VSS.n643 0.237342
R4835 VSS.n2177 VSS.n2176 0.237342
R4836 VSS.n2178 VSS.n2177 0.237342
R4837 VSS.n2178 VSS.n639 0.237342
R4838 VSS.n2184 VSS.n639 0.237342
R4839 VSS.n2185 VSS.n2184 0.237342
R4840 VSS.n2187 VSS.n2185 0.237342
R4841 VSS.n2187 VSS.n2186 0.237342
R4842 VSS.n2186 VSS.n635 0.237342
R4843 VSS.n2194 VSS.n635 0.237342
R4844 VSS.n2195 VSS.n2194 0.237342
R4845 VSS.n2196 VSS.n2195 0.237342
R4846 VSS.n2196 VSS.n629 0.237342
R4847 VSS.n588 VSS.n587 0.237342
R4848 VSS.n591 VSS.n588 0.237342
R4849 VSS.n592 VSS.n591 0.237342
R4850 VSS.n2334 VSS.n592 0.237342
R4851 VSS.n2334 VSS.n2333 0.237342
R4852 VSS.n2333 VSS.n2332 0.237342
R4853 VSS.n2332 VSS.n593 0.237342
R4854 VSS.n2326 VSS.n593 0.237342
R4855 VSS.n2326 VSS.n2325 0.237342
R4856 VSS.n2325 VSS.n2324 0.237342
R4857 VSS.n2324 VSS.n597 0.237342
R4858 VSS.n2318 VSS.n597 0.237342
R4859 VSS.n2318 VSS.n2317 0.237342
R4860 VSS.n2317 VSS.n2316 0.237342
R4861 VSS.n2316 VSS.n601 0.237342
R4862 VSS.n2310 VSS.n601 0.237342
R4863 VSS.n2310 VSS.n2309 0.237342
R4864 VSS.n2309 VSS.n2308 0.237342
R4865 VSS.n2308 VSS.n605 0.237342
R4866 VSS.n607 VSS.n605 0.237342
R4867 VSS.n2301 VSS.n607 0.237342
R4868 VSS.n517 VSS.n515 0.237342
R4869 VSS.n515 VSS.n472 0.237342
R4870 VSS.n2492 VSS.n472 0.237342
R4871 VSS.n2493 VSS.n2492 0.237342
R4872 VSS.n2494 VSS.n2493 0.237342
R4873 VSS.n2494 VSS.n468 0.237342
R4874 VSS.n2500 VSS.n468 0.237342
R4875 VSS.n2501 VSS.n2500 0.237342
R4876 VSS.n2502 VSS.n2501 0.237342
R4877 VSS.n2502 VSS.n464 0.237342
R4878 VSS.n2508 VSS.n464 0.237342
R4879 VSS.n2509 VSS.n2508 0.237342
R4880 VSS.n2510 VSS.n2509 0.237342
R4881 VSS.n2510 VSS.n460 0.237342
R4882 VSS.n2516 VSS.n460 0.237342
R4883 VSS.n2517 VSS.n2516 0.237342
R4884 VSS.n2523 VSS.n2517 0.237342
R4885 VSS.n2523 VSS.n2522 0.237342
R4886 VSS.n2522 VSS.n2521 0.237342
R4887 VSS.n2521 VSS.n2518 0.237342
R4888 VSS.n2518 VSS.n449 0.237342
R4889 VSS.n662 VSS.n64 0.237342
R4890 VSS.n668 VSS.n662 0.237342
R4891 VSS.n669 VSS.n668 0.237342
R4892 VSS.n682 VSS.n669 0.237342
R4893 VSS.n682 VSS.n681 0.237342
R4894 VSS.n681 VSS.n680 0.237342
R4895 VSS.n680 VSS.n677 0.237342
R4896 VSS.n677 VSS.n676 0.237342
R4897 VSS.n676 VSS.n673 0.237342
R4898 VSS.n673 VSS.n672 0.237342
R4899 VSS.n672 VSS.n670 0.237342
R4900 VSS.n670 VSS.n655 0.237342
R4901 VSS.n688 VSS.n655 0.237342
R4902 VSS.n689 VSS.n688 0.237342
R4903 VSS.n692 VSS.n689 0.237342
R4904 VSS.n693 VSS.n692 0.237342
R4905 VSS.n1673 VSS.n1672 0.237342
R4906 VSS.n1672 VSS.n1671 0.237342
R4907 VSS.n1671 VSS.n1574 0.237342
R4908 VSS.n1665 VSS.n1574 0.237342
R4909 VSS.n1665 VSS.n1664 0.237342
R4910 VSS.n1664 VSS.n1663 0.237342
R4911 VSS.n1663 VSS.n1629 0.237342
R4912 VSS.n1657 VSS.n1629 0.237342
R4913 VSS.n1655 VSS.n1654 0.237342
R4914 VSS.n1654 VSS.n1634 0.237342
R4915 VSS.n1648 VSS.n1634 0.237342
R4916 VSS.n1648 VSS.n1647 0.237342
R4917 VSS.n1647 VSS.n1646 0.237342
R4918 VSS.n1646 VSS.n1638 0.237342
R4919 VSS.n1640 VSS.n1638 0.237342
R4920 VSS.n1640 VSS.n809 0.237342
R4921 VSS.n1926 VSS.n809 0.237342
R4922 VSS.n1928 VSS.n804 0.237342
R4923 VSS.n1934 VSS.n804 0.237342
R4924 VSS.n1935 VSS.n1934 0.237342
R4925 VSS.n1936 VSS.n1935 0.237342
R4926 VSS.n1936 VSS.n800 0.237342
R4927 VSS.n1942 VSS.n800 0.237342
R4928 VSS.n1943 VSS.n1942 0.237342
R4929 VSS.n1946 VSS.n1943 0.237342
R4930 VSS.n1952 VSS.n796 0.237342
R4931 VSS.n1953 VSS.n1952 0.237342
R4932 VSS.n1954 VSS.n1953 0.237342
R4933 VSS.n1954 VSS.n792 0.237342
R4934 VSS.n1960 VSS.n792 0.237342
R4935 VSS.n1961 VSS.n1960 0.237342
R4936 VSS.n1962 VSS.n1961 0.237342
R4937 VSS.n1962 VSS.n788 0.237342
R4938 VSS.n1968 VSS.n788 0.237342
R4939 VSS.n2022 VSS.n1969 0.237342
R4940 VSS.n2016 VSS.n1969 0.237342
R4941 VSS.n2016 VSS.n2015 0.237342
R4942 VSS.n2015 VSS.n2014 0.237342
R4943 VSS.n2014 VSS.n1974 0.237342
R4944 VSS.n2008 VSS.n1974 0.237342
R4945 VSS.n2008 VSS.n2007 0.237342
R4946 VSS.n2007 VSS.n2006 0.237342
R4947 VSS.n2000 VSS.n1983 0.237342
R4948 VSS.n2000 VSS.n1999 0.237342
R4949 VSS.n1999 VSS.n1998 0.237342
R4950 VSS.n1998 VSS.n1984 0.237342
R4951 VSS.n1992 VSS.n1984 0.237342
R4952 VSS.n1992 VSS.n1991 0.237342
R4953 VSS.n1991 VSS.n1990 0.237342
R4954 VSS.n1990 VSS.n630 0.237342
R4955 VSS.n2203 VSS.n630 0.237342
R4956 VSS.n2205 VSS.n625 0.237342
R4957 VSS.n2211 VSS.n625 0.237342
R4958 VSS.n2212 VSS.n2211 0.237342
R4959 VSS.n2213 VSS.n2212 0.237342
R4960 VSS.n2213 VSS.n621 0.237342
R4961 VSS.n2219 VSS.n621 0.237342
R4962 VSS.n2220 VSS.n2219 0.237342
R4963 VSS.n2223 VSS.n2220 0.237342
R4964 VSS.n2229 VSS.n617 0.237342
R4965 VSS.n2230 VSS.n2229 0.237342
R4966 VSS.n2231 VSS.n2230 0.237342
R4967 VSS.n2231 VSS.n613 0.237342
R4968 VSS.n2237 VSS.n613 0.237342
R4969 VSS.n2238 VSS.n2237 0.237342
R4970 VSS.n2239 VSS.n2238 0.237342
R4971 VSS.n2239 VSS.n609 0.237342
R4972 VSS.n2245 VSS.n609 0.237342
R4973 VSS.n2299 VSS.n2246 0.237342
R4974 VSS.n2293 VSS.n2246 0.237342
R4975 VSS.n2293 VSS.n2292 0.237342
R4976 VSS.n2292 VSS.n2291 0.237342
R4977 VSS.n2291 VSS.n2251 0.237342
R4978 VSS.n2285 VSS.n2251 0.237342
R4979 VSS.n2285 VSS.n2284 0.237342
R4980 VSS.n2284 VSS.n2283 0.237342
R4981 VSS.n2277 VSS.n2260 0.237342
R4982 VSS.n2277 VSS.n2276 0.237342
R4983 VSS.n2276 VSS.n2275 0.237342
R4984 VSS.n2275 VSS.n2261 0.237342
R4985 VSS.n2269 VSS.n2261 0.237342
R4986 VSS.n2269 VSS.n2268 0.237342
R4987 VSS.n2268 VSS.n2267 0.237342
R4988 VSS.n2267 VSS.n450 0.237342
R4989 VSS.n2530 VSS.n450 0.237342
R4990 VSS.n2533 VSS.n2532 0.237342
R4991 VSS.n2533 VSS.n445 0.237342
R4992 VSS.n2539 VSS.n445 0.237342
R4993 VSS.n2540 VSS.n2539 0.237342
R4994 VSS.n2541 VSS.n2540 0.237342
R4995 VSS.n2541 VSS.n441 0.237342
R4996 VSS.n2547 VSS.n441 0.237342
R4997 VSS.n2548 VSS.n2547 0.237342
R4998 VSS.n2550 VSS.n436 0.237342
R4999 VSS.n2556 VSS.n436 0.237342
R5000 VSS.n2557 VSS.n2556 0.237342
R5001 VSS.n2558 VSS.n2557 0.237342
R5002 VSS.n2558 VSS.n432 0.237342
R5003 VSS.n2565 VSS.n432 0.237342
R5004 VSS.n2566 VSS.n2565 0.237342
R5005 VSS.n2567 VSS.n2566 0.237342
R5006 VSS.n2567 VSS.n424 0.237342
R5007 VSS.n2583 VSS.n420 0.237342
R5008 VSS.n2590 VSS.n420 0.237342
R5009 VSS.n2591 VSS.n2590 0.237342
R5010 VSS.n2592 VSS.n2591 0.237342
R5011 VSS.n2592 VSS.n415 0.237342
R5012 VSS.n2599 VSS.n415 0.237342
R5013 VSS.n2600 VSS.n2599 0.237342
R5014 VSS.n2602 VSS.n2600 0.237342
R5015 VSS.n2602 VSS.n2601 0.237342
R5016 VSS.n2609 VSS.n2608 0.237342
R5017 VSS.n2610 VSS.n2609 0.237342
R5018 VSS.n2610 VSS.n406 0.237342
R5019 VSS.n2616 VSS.n406 0.237342
R5020 VSS.n2617 VSS.n2616 0.237342
R5021 VSS.n2618 VSS.n2617 0.237342
R5022 VSS.n2618 VSS.n401 0.237342
R5023 VSS.n2654 VSS.n401 0.237342
R5024 VSS.n2658 VSS.n2656 0.237342
R5025 VSS.n2658 VSS.n2657 0.237342
R5026 VSS.n2657 VSS.n396 0.237342
R5027 VSS.n2665 VSS.n396 0.237342
R5028 VSS.n2666 VSS.n2665 0.237342
R5029 VSS.n2695 VSS.n2666 0.237342
R5030 VSS.n2695 VSS.n2694 0.237342
R5031 VSS.n2694 VSS.n2693 0.237342
R5032 VSS.n2693 VSS.n2667 0.237342
R5033 VSS.n2687 VSS.n2667 0.237342
R5034 VSS.n2687 VSS.n2686 0.237342
R5035 VSS.n2686 VSS.n2685 0.237342
R5036 VSS.n2685 VSS.n2671 0.237342
R5037 VSS.n2679 VSS.n2671 0.237342
R5038 VSS.n2679 VSS.n2678 0.237342
R5039 VSS.n2678 VSS.n2677 0.237342
R5040 VSS.n2677 VSS.n121 0.237342
R5041 VSS.n3241 VSS.n121 0.237342
R5042 VSS.n2402 VSS.n261 0.237342
R5043 VSS.n2408 VSS.n2402 0.237342
R5044 VSS.n2409 VSS.n2408 0.237342
R5045 VSS.n2444 VSS.n2409 0.237342
R5046 VSS.n2444 VSS.n2443 0.237342
R5047 VSS.n2443 VSS.n2442 0.237342
R5048 VSS.n2442 VSS.n2410 0.237342
R5049 VSS.n2436 VSS.n2410 0.237342
R5050 VSS.n2436 VSS.n2435 0.237342
R5051 VSS.n2435 VSS.n2434 0.237342
R5052 VSS.n2434 VSS.n2416 0.237342
R5053 VSS.n2420 VSS.n2416 0.237342
R5054 VSS.n2426 VSS.n2420 0.237342
R5055 VSS.n2426 VSS.n2425 0.237342
R5056 VSS.n2425 VSS.n2424 0.237342
R5057 VSS.n2424 VSS.n2421 0.237342
R5058 VSS.n2421 VSS.n427 0.237342
R5059 VSS.n2575 VSS.n427 0.237342
R5060 VSS.n2576 VSS.n2575 0.237342
R5061 VSS.n2576 VSS.n425 0.237342
R5062 VSS.n2581 VSS.n425 0.237342
R5063 VSS.n1782 VSS.n1781 0.237342
R5064 VSS.n1781 VSS.n1780 0.237342
R5065 VSS.n1780 VSS.n1733 0.237342
R5066 VSS.n1737 VSS.n1733 0.237342
R5067 VSS.n1773 VSS.n1737 0.237342
R5068 VSS.n1773 VSS.n1772 0.237342
R5069 VSS.n1772 VSS.n1771 0.237342
R5070 VSS.n1771 VSS.n1738 0.237342
R5071 VSS.n1765 VSS.n1738 0.237342
R5072 VSS.n1765 VSS.n1764 0.237342
R5073 VSS.n1764 VSS.n1763 0.237342
R5074 VSS.n1763 VSS.n1742 0.237342
R5075 VSS.n1757 VSS.n1742 0.237342
R5076 VSS.n1757 VSS.n1756 0.237342
R5077 VSS.n1756 VSS.n1755 0.237342
R5078 VSS.n1755 VSS.n1746 0.237342
R5079 VSS.n1749 VSS.n1746 0.237342
R5080 VSS.n1749 VSS.n1748 0.237342
R5081 VSS.n839 VSS.n836 0.237342
R5082 VSS.n881 VSS.n839 0.237342
R5083 VSS.n881 VSS.n880 0.237342
R5084 VSS.n880 VSS.n879 0.237342
R5085 VSS.n879 VSS.n840 0.237342
R5086 VSS.n873 VSS.n840 0.237342
R5087 VSS.n873 VSS.n872 0.237342
R5088 VSS.n872 VSS.n871 0.237342
R5089 VSS.n871 VSS.n844 0.237342
R5090 VSS.n865 VSS.n844 0.237342
R5091 VSS.n865 VSS.n864 0.237342
R5092 VSS.n864 VSS.n863 0.237342
R5093 VSS.n863 VSS.n848 0.237342
R5094 VSS.n857 VSS.n848 0.237342
R5095 VSS.n857 VSS.n856 0.237342
R5096 VSS.n856 VSS.n855 0.237342
R5097 VSS.n855 VSS.n852 0.237342
R5098 VSS.n852 VSS.n717 0.237342
R5099 VSS.n2069 VSS.n713 0.237342
R5100 VSS.n2070 VSS.n2069 0.237342
R5101 VSS.n2071 VSS.n2070 0.237342
R5102 VSS.n2071 VSS.n709 0.237342
R5103 VSS.n2077 VSS.n709 0.237342
R5104 VSS.n2078 VSS.n2077 0.237342
R5105 VSS.n2079 VSS.n2078 0.237342
R5106 VSS.n2079 VSS.n705 0.237342
R5107 VSS.n2085 VSS.n705 0.237342
R5108 VSS.n2086 VSS.n2085 0.237342
R5109 VSS.n2087 VSS.n2086 0.237342
R5110 VSS.n2087 VSS.n701 0.237342
R5111 VSS.n2093 VSS.n701 0.237342
R5112 VSS.n2094 VSS.n2093 0.237342
R5113 VSS.n2096 VSS.n2094 0.237342
R5114 VSS.n2096 VSS.n2095 0.237342
R5115 VSS.n2095 VSS.n698 0.237342
R5116 VSS.n698 VSS.n694 0.237342
R5117 VSS.n2154 VSS.n695 0.237342
R5118 VSS.n2148 VSS.n695 0.237342
R5119 VSS.n2148 VSS.n2147 0.237342
R5120 VSS.n2147 VSS.n2146 0.237342
R5121 VSS.n2146 VSS.n2107 0.237342
R5122 VSS.n2140 VSS.n2107 0.237342
R5123 VSS.n2140 VSS.n2139 0.237342
R5124 VSS.n2139 VSS.n2138 0.237342
R5125 VSS.n2138 VSS.n2111 0.237342
R5126 VSS.n2132 VSS.n2111 0.237342
R5127 VSS.n2132 VSS.n2131 0.237342
R5128 VSS.n2131 VSS.n2130 0.237342
R5129 VSS.n2130 VSS.n2115 0.237342
R5130 VSS.n2124 VSS.n2115 0.237342
R5131 VSS.n2124 VSS.n2123 0.237342
R5132 VSS.n2123 VSS.n2122 0.237342
R5133 VSS.n2122 VSS.n2119 0.237342
R5134 VSS.n2119 VSS.n538 0.237342
R5135 VSS.n2346 VSS.n534 0.237342
R5136 VSS.n2347 VSS.n2346 0.237342
R5137 VSS.n2348 VSS.n2347 0.237342
R5138 VSS.n2348 VSS.n530 0.237342
R5139 VSS.n2354 VSS.n530 0.237342
R5140 VSS.n2355 VSS.n2354 0.237342
R5141 VSS.n2356 VSS.n2355 0.237342
R5142 VSS.n2356 VSS.n526 0.237342
R5143 VSS.n2362 VSS.n526 0.237342
R5144 VSS.n2363 VSS.n2362 0.237342
R5145 VSS.n2364 VSS.n2363 0.237342
R5146 VSS.n2364 VSS.n522 0.237342
R5147 VSS.n2370 VSS.n522 0.237342
R5148 VSS.n2371 VSS.n2370 0.237342
R5149 VSS.n2373 VSS.n2371 0.237342
R5150 VSS.n2373 VSS.n2372 0.237342
R5151 VSS.n2372 VSS.n518 0.237342
R5152 VSS.n2380 VSS.n518 0.237342
R5153 VSS.n2484 VSS.n2381 0.237342
R5154 VSS.n2385 VSS.n2381 0.237342
R5155 VSS.n2477 VSS.n2385 0.237342
R5156 VSS.n2477 VSS.n2476 0.237342
R5157 VSS.n2476 VSS.n2475 0.237342
R5158 VSS.n2475 VSS.n2386 0.237342
R5159 VSS.n2469 VSS.n2386 0.237342
R5160 VSS.n2469 VSS.n2468 0.237342
R5161 VSS.n2468 VSS.n2467 0.237342
R5162 VSS.n2467 VSS.n2390 0.237342
R5163 VSS.n2461 VSS.n2390 0.237342
R5164 VSS.n2461 VSS.n2460 0.237342
R5165 VSS.n2460 VSS.n2459 0.237342
R5166 VSS.n2459 VSS.n2394 0.237342
R5167 VSS.n2453 VSS.n2394 0.237342
R5168 VSS.n2453 VSS.n2452 0.237342
R5169 VSS.n2452 VSS.n2451 0.237342
R5170 VSS.n2451 VSS.n262 0.237342
R5171 VSS.n2745 VSS.n263 0.237342
R5172 VSS.n2739 VSS.n263 0.237342
R5173 VSS.n2739 VSS.n2738 0.237342
R5174 VSS.n2738 VSS.n2737 0.237342
R5175 VSS.n2737 VSS.n267 0.237342
R5176 VSS.n269 VSS.n267 0.237342
R5177 VSS.n2730 VSS.n269 0.237342
R5178 VSS.n2730 VSS.n2729 0.237342
R5179 VSS.n2729 VSS.n2728 0.237342
R5180 VSS.n2728 VSS.n271 0.237342
R5181 VSS.n2722 VSS.n271 0.237342
R5182 VSS.n2722 VSS.n2721 0.237342
R5183 VSS.n2721 VSS.n2720 0.237342
R5184 VSS.n2720 VSS.n280 0.237342
R5185 VSS.n2714 VSS.n280 0.237342
R5186 VSS.n2714 VSS.n2713 0.237342
R5187 VSS.n2713 VSS.n2712 0.237342
R5188 VSS.n2712 VSS.n284 0.237342
R5189 VSS.n370 VSS.n369 0.237342
R5190 VSS.n370 VSS.n298 0.237342
R5191 VSS.n376 VSS.n298 0.237342
R5192 VSS.n377 VSS.n376 0.237342
R5193 VSS.n388 VSS.n377 0.237342
R5194 VSS.n388 VSS.n387 0.237342
R5195 VSS.n387 VSS.n386 0.237342
R5196 VSS.n386 VSS.n378 0.237342
R5197 VSS.n380 VSS.n378 0.237342
R5198 VSS.n380 VSS.n135 0.237342
R5199 VSS.n3219 VSS.n135 0.237342
R5200 VSS.n3219 VSS.n3218 0.237342
R5201 VSS.n3218 VSS.n3217 0.237342
R5202 VSS.n3217 VSS.n136 0.237342
R5203 VSS.n137 VSS.n136 0.237342
R5204 VSS.n3210 VSS.n137 0.237342
R5205 VSS.n3210 VSS.n3209 0.237342
R5206 VSS.n3209 VSS.n3208 0.237342
R5207 VSS.n733 VSS.n42 0.237342
R5208 VSS.n739 VSS.n733 0.237342
R5209 VSS.n740 VSS.n739 0.237342
R5210 VSS.n753 VSS.n740 0.237342
R5211 VSS.n753 VSS.n752 0.237342
R5212 VSS.n752 VSS.n751 0.237342
R5213 VSS.n751 VSS.n748 0.237342
R5214 VSS.n748 VSS.n747 0.237342
R5215 VSS.n747 VSS.n744 0.237342
R5216 VSS.n744 VSS.n743 0.237342
R5217 VSS.n743 VSS.n741 0.237342
R5218 VSS.n741 VSS.n726 0.237342
R5219 VSS.n759 VSS.n726 0.237342
R5220 VSS.n760 VSS.n759 0.237342
R5221 VSS.n763 VSS.n760 0.237342
R5222 VSS.n764 VSS.n763 0.237342
R5223 VSS.n1819 VSS.n1818 0.237342
R5224 VSS.n1834 VSS.n1819 0.237342
R5225 VSS.n1834 VSS.n1833 0.237342
R5226 VSS.n1833 VSS.n1832 0.237342
R5227 VSS.n1832 VSS.n1820 0.237342
R5228 VSS.n1826 VSS.n1820 0.237342
R5229 VSS.n1826 VSS.n1825 0.237342
R5230 VSS.n1825 VSS.n7 0.237342
R5231 VSS.n3424 VSS.n7 0.237342
R5232 VSS.n3422 VSS.n3421 0.237342
R5233 VSS.n3421 VSS.n10 0.237342
R5234 VSS.n3415 VSS.n10 0.237342
R5235 VSS.n3415 VSS.n3414 0.237342
R5236 VSS.n3414 VSS.n3413 0.237342
R5237 VSS.n3413 VSS.n15 0.237342
R5238 VSS.n3407 VSS.n15 0.237342
R5239 VSS.n3407 VSS.n3406 0.237342
R5240 VSS.n3404 VSS.n20 0.237342
R5241 VSS.n3398 VSS.n20 0.237342
R5242 VSS.n3398 VSS.n3397 0.237342
R5243 VSS.n3397 VSS.n3396 0.237342
R5244 VSS.n3396 VSS.n26 0.237342
R5245 VSS.n3390 VSS.n26 0.237342
R5246 VSS.n3390 VSS.n3389 0.237342
R5247 VSS.n3389 VSS.n3388 0.237342
R5248 VSS.n3388 VSS.n30 0.237342
R5249 VSS.n3382 VSS.n30 0.237342
R5250 VSS.n3382 VSS.n3381 0.237342
R5251 VSS.n3381 VSS.n3380 0.237342
R5252 VSS.n3380 VSS.n34 0.237342
R5253 VSS.n3374 VSS.n34 0.237342
R5254 VSS.n3374 VSS.n3373 0.237342
R5255 VSS.n3373 VSS.n3372 0.237342
R5256 VSS.n3372 VSS.n38 0.237342
R5257 VSS.n3366 VSS.n38 0.237342
R5258 VSS.n3364 VSS.n43 0.237342
R5259 VSS.n3358 VSS.n43 0.237342
R5260 VSS.n3358 VSS.n3357 0.237342
R5261 VSS.n3357 VSS.n3356 0.237342
R5262 VSS.n3356 VSS.n48 0.237342
R5263 VSS.n3350 VSS.n48 0.237342
R5264 VSS.n3350 VSS.n3349 0.237342
R5265 VSS.n3349 VSS.n3348 0.237342
R5266 VSS.n3348 VSS.n52 0.237342
R5267 VSS.n3342 VSS.n52 0.237342
R5268 VSS.n3342 VSS.n3341 0.237342
R5269 VSS.n3341 VSS.n3340 0.237342
R5270 VSS.n3340 VSS.n56 0.237342
R5271 VSS.n3334 VSS.n56 0.237342
R5272 VSS.n3334 VSS.n3333 0.237342
R5273 VSS.n3333 VSS.n3332 0.237342
R5274 VSS.n3332 VSS.n60 0.237342
R5275 VSS.n3326 VSS.n60 0.237342
R5276 VSS.n3324 VSS.n65 0.237342
R5277 VSS.n3318 VSS.n65 0.237342
R5278 VSS.n3318 VSS.n3317 0.237342
R5279 VSS.n3317 VSS.n3316 0.237342
R5280 VSS.n3316 VSS.n70 0.237342
R5281 VSS.n3310 VSS.n70 0.237342
R5282 VSS.n3310 VSS.n3309 0.237342
R5283 VSS.n3309 VSS.n3308 0.237342
R5284 VSS.n3308 VSS.n74 0.237342
R5285 VSS.n3302 VSS.n74 0.237342
R5286 VSS.n3302 VSS.n3301 0.237342
R5287 VSS.n3301 VSS.n3300 0.237342
R5288 VSS.n3300 VSS.n78 0.237342
R5289 VSS.n3294 VSS.n78 0.237342
R5290 VSS.n3294 VSS.n3293 0.237342
R5291 VSS.n3293 VSS.n3292 0.237342
R5292 VSS.n3292 VSS.n82 0.237342
R5293 VSS.n3286 VSS.n82 0.237342
R5294 VSS.n3284 VSS.n87 0.237342
R5295 VSS.n3278 VSS.n87 0.237342
R5296 VSS.n3278 VSS.n3277 0.237342
R5297 VSS.n3277 VSS.n3276 0.237342
R5298 VSS.n3276 VSS.n92 0.237342
R5299 VSS.n3270 VSS.n92 0.237342
R5300 VSS.n3270 VSS.n3269 0.237342
R5301 VSS.n3269 VSS.n3268 0.237342
R5302 VSS.n3268 VSS.n95 0.237342
R5303 VSS.n205 VSS.n95 0.237342
R5304 VSS.n206 VSS.n205 0.237342
R5305 VSS.n206 VSS.n202 0.237342
R5306 VSS.n212 VSS.n202 0.237342
R5307 VSS.n213 VSS.n212 0.237342
R5308 VSS.n215 VSS.n213 0.237342
R5309 VSS.n215 VSS.n214 0.237342
R5310 VSS.n214 VSS.n198 0.237342
R5311 VSS.n222 VSS.n198 0.237342
R5312 VSS.n2817 VSS.n2816 0.237342
R5313 VSS.n2816 VSS.n2815 0.237342
R5314 VSS.n2815 VSS.n224 0.237342
R5315 VSS.n2809 VSS.n224 0.237342
R5316 VSS.n2809 VSS.n2808 0.237342
R5317 VSS.n2808 VSS.n2807 0.237342
R5318 VSS.n2807 VSS.n228 0.237342
R5319 VSS.n2801 VSS.n228 0.237342
R5320 VSS.n2801 VSS.n2800 0.237342
R5321 VSS.n2800 VSS.n2799 0.237342
R5322 VSS.n2799 VSS.n232 0.237342
R5323 VSS.n2793 VSS.n232 0.237342
R5324 VSS.n2793 VSS.n2792 0.237342
R5325 VSS.n2792 VSS.n2791 0.237342
R5326 VSS.n2791 VSS.n236 0.237342
R5327 VSS.n2785 VSS.n236 0.237342
R5328 VSS.n2785 VSS.n2784 0.237342
R5329 VSS.n2784 VSS.n2783 0.237342
R5330 VSS.n2777 VSS.n2776 0.237342
R5331 VSS.n2776 VSS.n2775 0.237342
R5332 VSS.n2775 VSS.n162 0.237342
R5333 VSS.n3121 VSS.n162 0.237342
R5334 VSS.n3122 VSS.n3121 0.237342
R5335 VSS.n3123 VSS.n3122 0.237342
R5336 VSS.n3123 VSS.n160 0.237342
R5337 VSS.n3128 VSS.n160 0.237342
R5338 VSS.n3129 VSS.n3128 0.237342
R5339 VSS.n3130 VSS.n3129 0.237342
R5340 VSS.n3130 VSS.n158 0.237342
R5341 VSS.n158 VSS.n157 0.237342
R5342 VSS.n3137 VSS.n157 0.237342
R5343 VSS.n3138 VSS.n3137 0.237342
R5344 VSS.n3139 VSS.n3138 0.237342
R5345 VSS.n3139 VSS.n155 0.237342
R5346 VSS.n155 VSS.n154 0.237342
R5347 VSS.n3146 VSS.n154 0.237342
R5348 VSS.n3148 VSS.n151 0.237342
R5349 VSS.n3154 VSS.n151 0.237342
R5350 VSS.n3155 VSS.n3154 0.237342
R5351 VSS.n3156 VSS.n3155 0.237342
R5352 VSS.n3156 VSS.n149 0.237342
R5353 VSS.n3162 VSS.n149 0.237342
R5354 VSS.n3163 VSS.n3162 0.237342
R5355 VSS.n3164 VSS.n3163 0.237342
R5356 VSS.n3164 VSS.n147 0.237342
R5357 VSS.n3170 VSS.n147 0.237342
R5358 VSS.n3171 VSS.n3170 0.237342
R5359 VSS.n3172 VSS.n3171 0.237342
R5360 VSS.n3172 VSS.n145 0.237342
R5361 VSS.n3178 VSS.n145 0.237342
R5362 VSS.n3179 VSS.n3178 0.237342
R5363 VSS.n3180 VSS.n3179 0.237342
R5364 VSS.n3180 VSS.n143 0.237342
R5365 VSS.n3185 VSS.n143 0.237342
R5366 VSS.n1801 VSS.n904 0.235007
R5367 VSS.t108 VSS.n2878 0.233316
R5368 VSS.n1548 VSS.n1004 0.229053
R5369 VSS.n1154 VSS.n1153 0.226684
R5370 VSS.n1552 VSS.n897 0.226498
R5371 VSS.n1708 VSS.n938 0.223034
R5372 VSS.n1168 VSS.n1015 0.218395
R5373 VSS.n1119 VSS.n1063 0.218395
R5374 VSS.n3040 VSS.n106 0.217142
R5375 VSS.n1194 VSS.n1073 0.207737
R5376 VSS.n1152 VSS.n1123 0.207737
R5377 VSS.n1689 VSS.n1688 0.207623
R5378 VSS.n3423 VSS.n3422 0.204184
R5379 VSS.n1561 VSS.n906 0.1994
R5380 VSS.n3231 VSS.n3230 0.193093
R5381 VSS.n3230 VSS.n3229 0.193093
R5382 VSS.n3249 VSS.n3248 0.193093
R5383 VSS.n3248 VSS.n3247 0.193093
R5384 VSS.n1471 VSS.n1004 0.192342
R5385 VSS.n1473 VSS.n1472 0.189974
R5386 VSS.n1080 VSS.n1077 0.187417
R5387 VSS.n1118 VSS.n1117 0.186075
R5388 VSS.n991 VSS.n990 0.183582
R5389 VSS.n961 VSS.n926 0.183582
R5390 VSS.n1724 VSS.n927 0.183582
R5391 VSS.n1212 VSS.n1211 0.183187
R5392 VSS.n1796 VSS.n1795 0.181768
R5393 VSS.n974 VSS.n973 0.175877
R5394 VSS.n1082 VSS.n1075 0.1697
R5395 VSS.n1232 VSS.n1231 0.1661
R5396 VSS.n1229 VSS.n1227 0.1661
R5397 VSS.n3188 VSS.n3187 0.165427
R5398 VSS.n956 VSS.n955 0.163548
R5399 VSS.n2636 VSS.n2627 0.161553
R5400 VSS.n836 VSS.n833 0.161553
R5401 VSS.n765 VSS.n713 0.161553
R5402 VSS.n2155 VSS.n2154 0.161553
R5403 VSS.n586 VSS.n534 0.161553
R5404 VSS.n2485 VSS.n2484 0.161553
R5405 VSS.n2746 VSS.n2745 0.161553
R5406 VSS.n369 VSS.n368 0.161553
R5407 VSS.n1515 VSS.n1005 0.161553
R5408 VSS.n1617 VSS.n1573 0.161236
R5409 VSS.n1731 VSS.n1730 0.156415
R5410 VSS.n1656 VSS.n1655 0.150895
R5411 VSS.n1945 VSS.n796 0.150895
R5412 VSS.n1983 VSS.n1979 0.150895
R5413 VSS.n2222 VSS.n617 0.150895
R5414 VSS.n2260 VSS.n2256 0.150895
R5415 VSS.n2550 VSS.n2549 0.150895
R5416 VSS.n1469 VSS.n1246 0.148156
R5417 VSS.n1928 VSS.n1927 0.147342
R5418 VSS.n2023 VSS.n2022 0.147342
R5419 VSS.n2205 VSS.n2204 0.147342
R5420 VSS.n2300 VSS.n2299 0.147342
R5421 VSS.n2532 VSS.n2531 0.147342
R5422 VSS.n2583 VSS.n2582 0.147342
R5423 VSS.n2656 VSS.n2655 0.147342
R5424 VSS.n3405 VSS.n3404 0.147342
R5425 VSS.n3365 VSS.n3364 0.147342
R5426 VSS.n3325 VSS.n3324 0.147342
R5427 VSS.n3285 VSS.n3284 0.147342
R5428 VSS.n2817 VSS.n223 0.147342
R5429 VSS.n2777 VSS.n239 0.147342
R5430 VSS.n3148 VSS.n3147 0.147342
R5431 VSS.n1242 VSS.n1073 0.144974
R5432 VSS.n948 VSS.n947 0.141048
R5433 VSS.n1450 VSS.n1449 0.14
R5434 VSS.n1449 VSS.n1448 0.14
R5435 VSS.n1448 VSS.n1300 0.14
R5436 VSS.n1444 VSS.n1300 0.14
R5437 VSS.n1444 VSS.n1443 0.14
R5438 VSS.n1443 VSS.n1442 0.14
R5439 VSS.n1442 VSS.n1308 0.14
R5440 VSS.n1438 VSS.n1308 0.14
R5441 VSS.n1438 VSS.n1437 0.14
R5442 VSS.n1437 VSS.n1436 0.14
R5443 VSS.n1436 VSS.n1317 0.14
R5444 VSS.n1432 VSS.n1317 0.14
R5445 VSS.n1432 VSS.n1431 0.14
R5446 VSS.n1431 VSS.n1430 0.14
R5447 VSS.n1430 VSS.n1326 0.14
R5448 VSS.n1426 VSS.n1326 0.14
R5449 VSS.n1426 VSS.n1425 0.14
R5450 VSS.n1425 VSS.n103 0.14
R5451 VSS.n2608 VSS.n411 0.139053
R5452 VSS.n960 VSS.n959 0.13889
R5453 VSS.n984 VSS.n983 0.138582
R5454 VSS.n952 VSS.n951 0.138582
R5455 VSS.n1694 VSS.n1693 0.138582
R5456 VSS.n1812 VSS.n901 0.137401
R5457 VSS.n975 VSS.n974 0.137349
R5458 VSS.n1243 VSS.n1242 0.13667
R5459 VSS.n1554 VSS.n1553 0.132545
R5460 VSS.n1153 VSS.n1152 0.131947
R5461 VSS.n1603 VSS.n919 0.128528
R5462 VSS.n982 VSS.n981 0.128411
R5463 VSS.n1927 VSS.n1926 0.128395
R5464 VSS.n2023 VSS.n1968 0.128395
R5465 VSS.n2204 VSS.n2203 0.128395
R5466 VSS.n2300 VSS.n2245 0.128395
R5467 VSS.n2531 VSS.n2530 0.128395
R5468 VSS.n2582 VSS.n424 0.128395
R5469 VSS.n2655 VSS.n2654 0.128395
R5470 VSS.n3406 VSS.n3405 0.128395
R5471 VSS.n3366 VSS.n3365 0.128395
R5472 VSS.n3326 VSS.n3325 0.128395
R5473 VSS.n3286 VSS.n3285 0.128395
R5474 VSS.n223 VSS.n222 0.128395
R5475 VSS.n2783 VSS.n239 0.128395
R5476 VSS.n3147 VSS.n3146 0.128395
R5477 VSS.n1606 VSS.n919 0.125993
R5478 VSS.n1707 VSS.n1706 0.125
R5479 VSS.n955 VSS.n954 0.123479
R5480 VSS.n3189 VSS.n3188 0.120757
R5481 VSS.n1693 VSS.n1692 0.120089
R5482 VSS.n1782 VSS.n1732 0.118921
R5483 VSS.n1238 VSS.n1077 0.118667
R5484 VSS.n950 VSS.n949 0.117315
R5485 VSS.n1474 VSS.n1473 0.116553
R5486 VSS.n3191 VSS.n142 0.114565
R5487 VSS.n986 VSS.n985 0.114233
R5488 VSS.n1748 VSS.n833 0.114184
R5489 VSS.n765 VSS.n717 0.114184
R5490 VSS.n2155 VSS.n694 0.114184
R5491 VSS.n586 VSS.n538 0.114184
R5492 VSS.n2485 VSS.n2380 0.114184
R5493 VSS.n2746 VSS.n262 0.114184
R5494 VSS.n368 VSS.n284 0.114184
R5495 VSS.n1690 VSS.n1689 0.113925
R5496 VSS.n3261 VSS.n104 0.1085
R5497 VSS.n3195 VSS.n115 0.108076
R5498 VSS.n3242 VSS.n120 0.106292
R5499 VSS.n1673 VSS.n1573 0.104711
R5500 VSS.n1818 VSS.n896 0.104711
R5501 VSS.n958 VSS.n957 0.10437
R5502 VSS.n2655 VSS.n400 0.102342
R5503 VSS.n1927 VSS.n808 0.102342
R5504 VSS.n2024 VSS.n2023 0.102342
R5505 VSS.n2204 VSS.n629 0.102342
R5506 VSS.n2301 VSS.n2300 0.102342
R5507 VSS.n2531 VSS.n449 0.102342
R5508 VSS.n2582 VSS.n2581 0.102342
R5509 VSS.n368 VSS.n367 0.101158
R5510 VSS.n1879 VSS.n833 0.101158
R5511 VSS.n766 VSS.n765 0.101158
R5512 VSS.n2156 VSS.n2155 0.101158
R5513 VSS.n587 VSS.n586 0.101158
R5514 VSS.n2485 VSS.n517 0.101158
R5515 VSS.n2746 VSS.n261 0.101158
R5516 VSS.n2601 VSS.n411 0.0987895
R5517 VSS.n1731 VSS.n923 0.0981056
R5518 VSS.n1496 VSS.n1015 0.0952368
R5519 VSS.n1492 VSS.n1063 0.0952368
R5520 VSS.n3227 VSS.n3226 0.095011
R5521 VSS.n1238 VSS.n1237 0.0948615
R5522 VSS.n1697 VSS.n1696 0.0941986
R5523 VSS.n3234 VSS.n3233 0.0933571
R5524 VSS.n3235 VSS.n3234 0.0933571
R5525 VSS.n3237 VSS.n120 0.0933571
R5526 VSS.n3238 VSS.n3237 0.0933571
R5527 VSS.n3200 VSS.n3199 0.0933571
R5528 VSS.n3201 VSS.n3200 0.0933571
R5529 VSS.n3202 VSS.n3198 0.0933571
R5530 VSS.n3202 VSS.n3201 0.0933571
R5531 VSS.n3186 VSS.n108 0.0933571
R5532 VSS.n3254 VSS.n108 0.0933571
R5533 VSS.n947 VSS.n946 0.0905
R5534 VSS.n2823 VSS.n2822 0.0895206
R5535 VSS.n3038 VSS.n106 0.0874537
R5536 VSS.n1657 VSS.n1656 0.0869474
R5537 VSS.n1946 VSS.n1945 0.0869474
R5538 VSS.n2006 VSS.n1979 0.0869474
R5539 VSS.n2223 VSS.n2222 0.0869474
R5540 VSS.n2283 VSS.n2256 0.0869474
R5541 VSS.n2549 VSS.n2548 0.0869474
R5542 VSS.n3405 VSS.n19 0.0833947
R5543 VSS.n3147 VSS.n153 0.0833947
R5544 VSS.n246 VSS.n239 0.0833947
R5545 VSS.n485 VSS.n223 0.0833947
R5546 VSS.n3285 VSS.n86 0.0833947
R5547 VSS.n3325 VSS.n64 0.0833947
R5548 VSS.n3365 VSS.n42 0.0833947
R5549 VSS VSS.n3430 0.0832564
R5550 VSS.n1472 VSS.n1471 0.08159
R5551 VSS.n988 VSS.n987 0.0797123
R5552 VSS.n1239 VSS.n1238 0.0772371
R5553 VSS.n1709 VSS.n937 0.0755346
R5554 VSS.n1227 VSS.n1226 0.0743
R5555 VSS.n1226 VSS.n1208 0.0743
R5556 VSS.n1557 VSS.n965 0.0743
R5557 VSS.n1558 VSS.n1557 0.0743
R5558 VSS.n1797 VSS.n1796 0.0727535
R5559 VSS.n971 VSS.n938 0.0695411
R5560 VSS.n959 VSS.n958 0.0692329
R5561 VSS.n1560 VSS.n1559 0.0689
R5562 VSS.n1223 VSS.n1222 0.0680325
R5563 VSS.n1224 VSS.n1223 0.0680325
R5564 VSS.n1081 VSS.n1080 0.0680325
R5565 VSS.n1112 VSS.n1081 0.0680325
R5566 VSS.n3189 VSS.n139 0.0626638
R5567 VSS.n1453 VSS.n1452 0.0626562
R5568 VSS.n954 VSS.n953 0.060911
R5569 VSS.n989 VSS.n988 0.0596781
R5570 VSS.n946 VSS.n939 0.0596781
R5571 VSS.n987 VSS.n986 0.0593699
R5572 VSS.n973 VSS.n972 0.0584452
R5573 VSS.n977 VSS.n976 0.0584452
R5574 VSS.n980 VSS.n979 0.0584452
R5575 VSS.n990 VSS.n989 0.0584452
R5576 VSS.n953 VSS.n952 0.0584452
R5577 VSS.n961 VSS.n960 0.0584452
R5578 VSS.n1688 VSS.n927 0.0584452
R5579 VSS.n3243 VSS.n3242 0.0576584
R5580 VSS.n3429 VSS.n3 0.0561818
R5581 VSS.n978 VSS.n977 0.0559795
R5582 VSS.n981 VSS.n980 0.0559795
R5583 VSS.n1696 VSS.n1695 0.0559795
R5584 VSS.n1722 VSS.n1721 0.0559198
R5585 VSS.n3196 VSS.n3194 0.0519837
R5586 VSS.n1704 VSS.n1703 0.0517977
R5587 VSS.n1703 VSS.n1702 0.0517977
R5588 VSS.n1702 VSS.n1701 0.0517977
R5589 VSS.n1701 VSS.n931 0.0517977
R5590 VSS.n1718 VSS.n1717 0.0517977
R5591 VSS.n1720 VSS.n1719 0.0517977
R5592 VSS.n1721 VSS.n1720 0.0517977
R5593 VSS.n1716 VSS.n931 0.0513397
R5594 VSS.n1473 VSS.n1004 0.0490526
R5595 VSS.n3426 VSS.n3425 0.0480786
R5596 VSS.n1214 VSS.n1213 0.0470589
R5597 VSS.n1221 VSS.n1220 0.0470589
R5598 VSS.n1218 VSS.n1217 0.0470589
R5599 VSS.n1217 VSS.n1216 0.0470589
R5600 VSS.n1216 VSS.n1215 0.0470589
R5601 VSS.n1215 VSS.n966 0.0470589
R5602 VSS.n1875 VSS.n833 0.0466842
R5603 VSS.n368 VSS.n302 0.0466842
R5604 VSS.n2747 VSS.n2746 0.0466842
R5605 VSS.n2486 VSS.n2485 0.0466842
R5606 VSS.n586 VSS.n585 0.0466842
R5607 VSS.n2155 VSS.n693 0.0466842
R5608 VSS.n765 VSS.n764 0.0466842
R5609 VSS.n3258 VSS.n3257 0.0461627
R5610 VSS.n1213 VSS.n1212 0.0459157
R5611 VSS.n1222 VSS.n1214 0.0438372
R5612 VSS.n1219 VSS.n992 0.0438333
R5613 VSS.n1210 VSS.n992 0.0438333
R5614 VSS.n1716 VSS.n1715 0.0438333
R5615 VSS.n1715 VSS.n1714 0.0438333
R5616 VSS.n1470 VSS.n1469 0.0423279
R5617 VSS.n1293 VSS.n1292 0.035375
R5618 VSS.n1452 VSS.n1296 0.035375
R5619 VSS.n1301 VSS.n1296 0.035375
R5620 VSS.n1303 VSS.n1301 0.035375
R5621 VSS.n1305 VSS.n1303 0.035375
R5622 VSS.n1309 VSS.n1305 0.035375
R5623 VSS.n1310 VSS.n1309 0.035375
R5624 VSS.n1312 VSS.n1310 0.035375
R5625 VSS.n1314 VSS.n1312 0.035375
R5626 VSS.n1318 VSS.n1314 0.035375
R5627 VSS.n1319 VSS.n1318 0.035375
R5628 VSS.n1321 VSS.n1319 0.035375
R5629 VSS.n1323 VSS.n1321 0.035375
R5630 VSS.n1327 VSS.n1323 0.035375
R5631 VSS.n1328 VSS.n1327 0.035375
R5632 VSS.n1330 VSS.n1328 0.035375
R5633 VSS.n1332 VSS.n1330 0.035375
R5634 VSS.n3424 VSS.n3423 0.0336579
R5635 VSS.n1711 VSS.n932 0.0318766
R5636 VSS.t108 VSS.n3041 0.0317616
R5637 VSS.n3226 VSS.n127 0.0317469
R5638 VSS.n1726 VSS.n1725 0.0314524
R5639 VSS.n1726 VSS.n912 0.0314524
R5640 VSS.n1706 VSS.n932 0.0314524
R5641 VSS.n3011 VSS.n3010 0.0303125
R5642 VSS.n3011 VSS.n2890 0.0303125
R5643 VSS.n3015 VSS.n2890 0.0303125
R5644 VSS.n3016 VSS.n3015 0.0303125
R5645 VSS.n3017 VSS.n3016 0.0303125
R5646 VSS.n3017 VSS.n2888 0.0303125
R5647 VSS.n3021 VSS.n2888 0.0303125
R5648 VSS.n3022 VSS.n3021 0.0303125
R5649 VSS.n3023 VSS.n3022 0.0303125
R5650 VSS.n3023 VSS.n2886 0.0303125
R5651 VSS.n3027 VSS.n2886 0.0303125
R5652 VSS.n3028 VSS.n3027 0.0303125
R5653 VSS.n3029 VSS.n3028 0.0303125
R5654 VSS.n3029 VSS.n2884 0.0303125
R5655 VSS.n3033 VSS.n2884 0.0303125
R5656 VSS.n3034 VSS.n3033 0.0303125
R5657 VSS.n3035 VSS.n3034 0.0303125
R5658 VSS.n3035 VSS.n2882 0.0303125
R5659 VSS.n3039 VSS.n2882 0.0303125
R5660 VSS.n3040 VSS.n3039 0.0303125
R5661 VSS.n3012 VSS.n2891 0.0303125
R5662 VSS.n3013 VSS.n3012 0.0303125
R5663 VSS.n3014 VSS.n3013 0.0303125
R5664 VSS.n3014 VSS.n2889 0.0303125
R5665 VSS.n3018 VSS.n2889 0.0303125
R5666 VSS.n3019 VSS.n3018 0.0303125
R5667 VSS.n3020 VSS.n3019 0.0303125
R5668 VSS.n3020 VSS.n2887 0.0303125
R5669 VSS.n3024 VSS.n2887 0.0303125
R5670 VSS.n3025 VSS.n3024 0.0303125
R5671 VSS.n3026 VSS.n3025 0.0303125
R5672 VSS.n3026 VSS.n2885 0.0303125
R5673 VSS.n3030 VSS.n2885 0.0303125
R5674 VSS.n3031 VSS.n3030 0.0303125
R5675 VSS.n3032 VSS.n3031 0.0303125
R5676 VSS.n3032 VSS.n2883 0.0303125
R5677 VSS.n3036 VSS.n2883 0.0303125
R5678 VSS.n3037 VSS.n3036 0.0303125
R5679 VSS.n3038 VSS.n3037 0.0303125
R5680 VSS.n951 VSS.n950 0.030089
R5681 VSS.n1237 VSS.n936 0.0300285
R5682 VSS.n3041 VSS.n3040 0.0299118
R5683 VSS.n2637 VSS.n2636 0.0289211
R5684 VSS.n1212 VSS.n937 0.028664
R5685 VSS.n1336 VSS.n1298 0.0284
R5686 VSS.n1336 VSS.n1302 0.0284
R5687 VSS.n1304 VSS.n1302 0.0284
R5688 VSS.n1306 VSS.n1304 0.0284
R5689 VSS.n1341 VSS.n1306 0.0284
R5690 VSS.n1341 VSS.n1311 0.0284
R5691 VSS.n1313 VSS.n1311 0.0284
R5692 VSS.n1315 VSS.n1313 0.0284
R5693 VSS.n1346 VSS.n1315 0.0284
R5694 VSS.n1346 VSS.n1320 0.0284
R5695 VSS.n1322 VSS.n1320 0.0284
R5696 VSS.n1324 VSS.n1322 0.0284
R5697 VSS.n1350 VSS.n1324 0.0284
R5698 VSS.n1350 VSS.n1329 0.0284
R5699 VSS.n1331 VSS.n1329 0.0284
R5700 VSS.n1333 VSS.n1331 0.0284
R5701 VSS.n1423 VSS.n1333 0.0284
R5702 VSS.n1423 VSS.n1422 0.0284
R5703 VSS.n1451 VSS.n1299 0.0284
R5704 VSS.n1447 VSS.n1299 0.0284
R5705 VSS.n1447 VSS.n1446 0.0284
R5706 VSS.n1446 VSS.n1445 0.0284
R5707 VSS.n1445 VSS.n1307 0.0284
R5708 VSS.n1441 VSS.n1307 0.0284
R5709 VSS.n1441 VSS.n1440 0.0284
R5710 VSS.n1440 VSS.n1439 0.0284
R5711 VSS.n1439 VSS.n1316 0.0284
R5712 VSS.n1435 VSS.n1316 0.0284
R5713 VSS.n1435 VSS.n1434 0.0284
R5714 VSS.n1434 VSS.n1433 0.0284
R5715 VSS.n1433 VSS.n1325 0.0284
R5716 VSS.n1429 VSS.n1325 0.0284
R5717 VSS.n1429 VSS.n1428 0.0284
R5718 VSS.n1428 VSS.n1427 0.0284
R5719 VSS.n1427 VSS.n1424 0.0284
R5720 VSS.n1219 VSS.n1218 0.0279365
R5721 VSS.n3008 VSS.n3005 0.0274686
R5722 VSS.n1240 VSS.n1239 0.02642
R5723 VSS.n1243 VSS.n1072 0.0258274
R5724 VSS.n979 VSS.n978 0.0251575
R5725 VSS.n985 VSS.n984 0.0248493
R5726 VSS.n3245 VSS.n3244 0.0245741
R5727 VSS.n3246 VSS.n3245 0.0245741
R5728 VSS.n1373 VSS.n1298 0.0239
R5729 VSS.n1451 VSS.n1297 0.0239
R5730 VSS.n926 VSS.n907 0.023
R5731 VSS.n3259 VSS.n106 0.0229864
R5732 VSS.n1719 VSS.n1718 0.0220267
R5733 VSS.n1723 VSS.n1722 0.0220267
R5734 VSS.n1338 VSS.n1337 0.0219615
R5735 VSS.n1339 VSS.n1338 0.0219615
R5736 VSS.n1340 VSS.n1339 0.0219615
R5737 VSS.n1342 VSS.n1340 0.0219615
R5738 VSS.n1343 VSS.n1342 0.0219615
R5739 VSS.n1344 VSS.n1343 0.0219615
R5740 VSS.n1345 VSS.n1344 0.0219615
R5741 VSS.t43 VSS.n1345 0.0219615
R5742 VSS.t43 VSS.n1354 0.0219615
R5743 VSS.n1354 VSS.n1353 0.0219615
R5744 VSS.n1353 VSS.n1352 0.0219615
R5745 VSS.n1352 VSS.n1351 0.0219615
R5746 VSS.n1351 VSS.n1349 0.0219615
R5747 VSS.n1349 VSS.n1348 0.0219615
R5748 VSS.n1348 VSS.n1347 0.0219615
R5749 VSS.n1347 VSS.n1335 0.0219615
R5750 VSS.n1420 VSS.n1335 0.0219615
R5751 VSS.n1288 VSS.n9 0.0215938
R5752 VSS.n1554 VSS.n966 0.0200381
R5753 VSS.n2826 VSS.n185 0.0199425
R5754 VSS.n3112 VSS.n185 0.0199425
R5755 VSS.n3112 VSS.n186 0.0199425
R5756 VSS.n3108 VSS.n186 0.0199425
R5757 VSS.n3108 VSS.n2828 0.0199425
R5758 VSS.n2832 VSS.n2828 0.0199425
R5759 VSS.n3100 VSS.n2832 0.0199425
R5760 VSS.n3100 VSS.n2833 0.0199425
R5761 VSS.n3096 VSS.n2833 0.0199425
R5762 VSS.n3096 VSS.n2837 0.0199425
R5763 VSS.n3090 VSS.n2837 0.0199425
R5764 VSS.n3090 VSS.n2840 0.0199425
R5765 VSS.n3086 VSS.n2840 0.0199425
R5766 VSS.n3086 VSS.n2843 0.0199425
R5767 VSS.n3080 VSS.n2843 0.0199425
R5768 VSS.n3080 VSS.n2847 0.0199425
R5769 VSS.n3076 VSS.n2847 0.0199425
R5770 VSS.n3076 VSS.n2848 0.0199425
R5771 VSS.n3070 VSS.n2848 0.0199425
R5772 VSS.n3070 VSS.n2853 0.0199425
R5773 VSS.n3066 VSS.n2853 0.0199425
R5774 VSS.n3066 VSS.n2856 0.0199425
R5775 VSS.n2858 VSS.n2856 0.0199425
R5776 VSS.n2861 VSS.n2858 0.0199425
R5777 VSS.n3056 VSS.n2861 0.0199425
R5778 VSS.n3056 VSS.n2862 0.0199425
R5779 VSS.n3052 VSS.n2862 0.0199425
R5780 VSS.n3052 VSS.n2865 0.0199425
R5781 VSS.n3046 VSS.n2865 0.0199425
R5782 VSS.n3046 VSS.n2868 0.0199425
R5783 VSS.n2922 VSS.n2868 0.0199425
R5784 VSS.n2922 VSS.n2921 0.0199425
R5785 VSS.n2921 VSS.n2917 0.0199425
R5786 VSS.n2933 VSS.n2917 0.0199425
R5787 VSS.n2933 VSS.n2915 0.0199425
R5788 VSS.n2937 VSS.n2915 0.0199425
R5789 VSS.n2938 VSS.n2937 0.0199425
R5790 VSS.n2938 VSS.n2912 0.0199425
R5791 VSS.n2945 VSS.n2912 0.0199425
R5792 VSS.n2945 VSS.n2911 0.0199425
R5793 VSS.n2950 VSS.n2911 0.0199425
R5794 VSS.n2950 VSS.n2908 0.0199425
R5795 VSS.n2956 VSS.n2908 0.0199425
R5796 VSS.n2957 VSS.n2956 0.0199425
R5797 VSS.n2963 VSS.n2957 0.0199425
R5798 VSS.n2963 VSS.n2958 0.0199425
R5799 VSS.n2958 VSS.n2905 0.0199425
R5800 VSS.n2905 VSS.n2902 0.0199425
R5801 VSS.n2974 VSS.n2902 0.0199425
R5802 VSS.n2975 VSS.n2974 0.0199425
R5803 VSS.n2976 VSS.n2975 0.0199425
R5804 VSS.n2976 VSS.n2899 0.0199425
R5805 VSS.n2983 VSS.n2899 0.0199425
R5806 VSS.n2983 VSS.n2897 0.0199425
R5807 VSS.n2987 VSS.n2897 0.0199425
R5808 VSS.n2987 VSS.n2894 0.0199425
R5809 VSS.n2994 VSS.n2894 0.0199425
R5810 VSS.n2995 VSS.n2994 0.0199425
R5811 VSS.n3000 VSS.n2995 0.0199425
R5812 VSS.n3000 VSS.n2996 0.0199425
R5813 VSS.n2996 VSS.n2881 0.0199425
R5814 VSS.n2825 VSS.n183 0.0199425
R5815 VSS.n3113 VSS.n183 0.0199425
R5816 VSS.n3113 VSS.n184 0.0199425
R5817 VSS.n3107 VSS.n184 0.0199425
R5818 VSS.n3107 VSS.n3105 0.0199425
R5819 VSS.n3105 VSS.n2829 0.0199425
R5820 VSS.n3101 VSS.n2829 0.0199425
R5821 VSS.n3101 VSS.n2831 0.0199425
R5822 VSS.n3095 VSS.n2831 0.0199425
R5823 VSS.n3095 VSS.n2838 0.0199425
R5824 VSS.n3091 VSS.n2838 0.0199425
R5825 VSS.n3091 VSS.n2839 0.0199425
R5826 VSS.n3085 VSS.n2839 0.0199425
R5827 VSS.n3085 VSS.n2844 0.0199425
R5828 VSS.n3081 VSS.n2844 0.0199425
R5829 VSS.n3081 VSS.n2846 0.0199425
R5830 VSS.n3075 VSS.n2846 0.0199425
R5831 VSS.n3075 VSS.n2849 0.0199425
R5832 VSS.n3071 VSS.n2849 0.0199425
R5833 VSS.n3071 VSS.n2852 0.0199425
R5834 VSS.n3065 VSS.n2852 0.0199425
R5835 VSS.n3065 VSS.n3062 0.0199425
R5836 VSS.n3062 VSS.n3061 0.0199425
R5837 VSS.n3061 VSS.n2857 0.0199425
R5838 VSS.n3057 VSS.n2857 0.0199425
R5839 VSS.n3057 VSS.n2860 0.0199425
R5840 VSS.n3051 VSS.n2860 0.0199425
R5841 VSS.n3051 VSS.n2866 0.0199425
R5842 VSS.n3047 VSS.n2866 0.0199425
R5843 VSS.n3047 VSS.n2867 0.0199425
R5844 VSS.n2923 VSS.n2867 0.0199425
R5845 VSS.n2923 VSS.n2918 0.0199425
R5846 VSS.n2927 VSS.n2918 0.0199425
R5847 VSS.n2932 VSS.n2927 0.0199425
R5848 VSS.n2932 VSS.n2928 0.0199425
R5849 VSS.n2928 VSS.n2914 0.0199425
R5850 VSS.n2939 VSS.n2914 0.0199425
R5851 VSS.n2939 VSS.n2913 0.0199425
R5852 VSS.n2944 VSS.n2913 0.0199425
R5853 VSS.n2944 VSS.n2910 0.0199425
R5854 VSS.n2951 VSS.n2910 0.0199425
R5855 VSS.n2951 VSS.n2909 0.0199425
R5856 VSS.n2955 VSS.n2909 0.0199425
R5857 VSS.n2955 VSS.n2907 0.0199425
R5858 VSS.n2964 VSS.n2907 0.0199425
R5859 VSS.n2964 VSS.n2904 0.0199425
R5860 VSS.n2968 VSS.n2904 0.0199425
R5861 VSS.n2969 VSS.n2968 0.0199425
R5862 VSS.n2973 VSS.n2969 0.0199425
R5863 VSS.n2973 VSS.n2901 0.0199425
R5864 VSS.n2977 VSS.n2901 0.0199425
R5865 VSS.n2977 VSS.n2900 0.0199425
R5866 VSS.n2982 VSS.n2900 0.0199425
R5867 VSS.n2982 VSS.n2896 0.0199425
R5868 VSS.n2988 VSS.n2896 0.0199425
R5869 VSS.n2988 VSS.n2895 0.0199425
R5870 VSS.n2993 VSS.n2895 0.0199425
R5871 VSS.n2993 VSS.n2893 0.0199425
R5872 VSS.n3001 VSS.n2893 0.0199425
R5873 VSS.n3001 VSS.n2892 0.0199425
R5874 VSS.n3005 VSS.n2892 0.0199425
R5875 VSS.n1469 VSS.n1468 0.0198648
R5876 VSS.n1220 VSS.n1219 0.0196224
R5877 VSS.n1797 VSS.n904 0.0195141
R5878 VSS.t43 VSS.n1337 0.0191923
R5879 VSS.n1470 VSS.n1244 0.0189426
R5880 VSS.n3263 VSS.n3262 0.0188746
R5881 VSS.n3264 VSS.n3263 0.0188746
R5882 VSS.n1370 VSS.n1369 0.0183702
R5883 VSS.n1369 VSS.n1290 0.0183702
R5884 VSS.n1368 VSS.n1366 0.0183702
R5885 VSS.n1366 VSS.n1289 0.0183702
R5886 VSS.n1365 VSS.n1288 0.0183702
R5887 VSS.n1453 VSS.n1294 0.0183702
R5888 VSS.n1370 VSS.n1246 0.0183702
R5889 VSS.n1368 VSS.n1367 0.0183702
R5890 VSS.n1365 VSS.n1364 0.0183702
R5891 VSS.n1294 VSS.n1293 0.0183702
R5892 VSS.n1367 VSS.n1290 0.0183702
R5893 VSS.n1364 VSS.n1289 0.0183702
R5894 VSS.n2824 VSS.n181 0.0176692
R5895 VSS.n3114 VSS.n182 0.0176692
R5896 VSS.n3106 VSS.n182 0.0176692
R5897 VSS.n3104 VSS.n3103 0.0176692
R5898 VSS.n3103 VSS.n3102 0.0176692
R5899 VSS.n3102 VSS.n2830 0.0176692
R5900 VSS.n3094 VSS.n3093 0.0176692
R5901 VSS.n3093 VSS.n3092 0.0176692
R5902 VSS.n3084 VSS.n2845 0.0176692
R5903 VSS.n3084 VSS.n3083 0.0176692
R5904 VSS.n3083 VSS.n3082 0.0176692
R5905 VSS.n3074 VSS.n2850 0.0176692
R5906 VSS.n3074 VSS.n3073 0.0176692
R5907 VSS.n3073 VSS.n3072 0.0176692
R5908 VSS.n3072 VSS.n2851 0.0176692
R5909 VSS.n3064 VSS.n2851 0.0176692
R5910 VSS.n3064 VSS.n3063 0.0176692
R5911 VSS.n3060 VSS.n3059 0.0176692
R5912 VSS.n3059 VSS.n3058 0.0176692
R5913 VSS.n3058 VSS.n2859 0.0176692
R5914 VSS.n3050 VSS.n3049 0.0176692
R5915 VSS.n3049 VSS.n3048 0.0176692
R5916 VSS.n2924 VSS.n2919 0.0176692
R5917 VSS.n2925 VSS.n2924 0.0176692
R5918 VSS.n2926 VSS.n2925 0.0176692
R5919 VSS.n2931 VSS.n2930 0.0176692
R5920 VSS.n2930 VSS.n2929 0.0176692
R5921 VSS.n2941 VSS.n2940 0.0176692
R5922 VSS.n2943 VSS.n2941 0.0176692
R5923 VSS.n2943 VSS.n2942 0.0176692
R5924 VSS.n2953 VSS.n2952 0.0176692
R5925 VSS.n2954 VSS.n2953 0.0176692
R5926 VSS.n2965 VSS.n2906 0.0176692
R5927 VSS.n2966 VSS.n2965 0.0176692
R5928 VSS.n2967 VSS.n2966 0.0176692
R5929 VSS.n2972 VSS.n2970 0.0176692
R5930 VSS.n2972 VSS.n2971 0.0176692
R5931 VSS.n2979 VSS.n2978 0.0176692
R5932 VSS.n2981 VSS.n2979 0.0176692
R5933 VSS.n2981 VSS.n2980 0.0176692
R5934 VSS.n2990 VSS.n2989 0.0176692
R5935 VSS.n2992 VSS.n2990 0.0176692
R5936 VSS.n2992 VSS.n2991 0.0176692
R5937 VSS.n3003 VSS.n3002 0.0176692
R5938 VSS.n3004 VSS.n3003 0.0176692
R5939 VSS.n2971 VSS.n171 0.0173923
R5940 VSS.n3009 VSS.n3008 0.0171202
R5941 VSS.n3092 VSS.n166 0.0168385
R5942 VSS.n2827 VSS.n187 0.0165807
R5943 VSS.n3111 VSS.n187 0.0165807
R5944 VSS.n3111 VSS.n3110 0.0165807
R5945 VSS.n3110 VSS.n3109 0.0165807
R5946 VSS.n2835 VSS.n2834 0.0165807
R5947 VSS.n3099 VSS.n2835 0.0165807
R5948 VSS.n3099 VSS.n3098 0.0165807
R5949 VSS.n3098 VSS.n3097 0.0165807
R5950 VSS.n3097 VSS.n2836 0.0165807
R5951 VSS.n3089 VSS.n3088 0.0165807
R5952 VSS.n3088 VSS.n3087 0.0165807
R5953 VSS.n3087 VSS.n2842 0.0165807
R5954 VSS.n3079 VSS.n2842 0.0165807
R5955 VSS.n3079 VSS.n3078 0.0165807
R5956 VSS.n3078 VSS.n3077 0.0165807
R5957 VSS.n3069 VSS.n2854 0.0165807
R5958 VSS.n3069 VSS.n3068 0.0165807
R5959 VSS.n3068 VSS.n3067 0.0165807
R5960 VSS.n3067 VSS.n2855 0.0165807
R5961 VSS.n2870 VSS.n2855 0.0165807
R5962 VSS.n3055 VSS.n2863 0.0165807
R5963 VSS.n3055 VSS.n3054 0.0165807
R5964 VSS.n3054 VSS.n3053 0.0165807
R5965 VSS.n3053 VSS.n2864 0.0165807
R5966 VSS.n3045 VSS.n2864 0.0165807
R5967 VSS.n3045 VSS.n3044 0.0165807
R5968 VSS.n2920 VSS.n2869 0.0165807
R5969 VSS.n2920 VSS.n2916 0.0165807
R5970 VSS.n2934 VSS.n2916 0.0165807
R5971 VSS.n2935 VSS.n2934 0.0165807
R5972 VSS.n2936 VSS.n2935 0.0165807
R5973 VSS.n2936 VSS.n2872 0.0165807
R5974 VSS.n2946 VSS.n2873 0.0165807
R5975 VSS.n2947 VSS.n2946 0.0165807
R5976 VSS.n2949 VSS.n2947 0.0165807
R5977 VSS.n2949 VSS.n2948 0.0165807
R5978 VSS.n2948 VSS.n2874 0.0165807
R5979 VSS.n2962 VSS.n2875 0.0165807
R5980 VSS.n2962 VSS.n2961 0.0165807
R5981 VSS.n2961 VSS.n2960 0.0165807
R5982 VSS.n2960 VSS.n2959 0.0165807
R5983 VSS.n2959 VSS.n2903 0.0165807
R5984 VSS.n2903 VSS.n2876 0.0165807
R5985 VSS.n2898 VSS.n2877 0.0165807
R5986 VSS.n2984 VSS.n2898 0.0165807
R5987 VSS.n2985 VSS.n2984 0.0165807
R5988 VSS.n2986 VSS.n2985 0.0165807
R5989 VSS.n2986 VSS.n2879 0.0165807
R5990 VSS.n2997 VSS.n2880 0.0165807
R5991 VSS.n2999 VSS.n2997 0.0165807
R5992 VSS.n2999 VSS.n2998 0.0165807
R5993 VSS.n2998 VSS.n2878 0.0165807
R5994 VSS.n3002 VSS.n172 0.0162846
R5995 VSS.n3430 VSS.n3429 0.0159762
R5996 VSS.n3429 VSS.n3428 0.0159762
R5997 VSS.n3260 VSS.n105 0.0158232
R5998 VSS.n2834 VSS.t209 0.0158026
R5999 VSS.t108 VSS.n2879 0.0158026
R6000 VSS.n2954 VSS.n170 0.0157308
R6001 VSS.n3244 VSS.n116 0.0154357
R6002 VSS.n3106 VSS.n165 0.0151769
R6003 VSS.n3050 VSS.n178 0.0151769
R6004 VSS.n3007 VSS.n3006 0.0151769
R6005 VSS.n139 VSS.n127 0.0151333
R6006 VSS.n1421 VSS.n1334 0.0149713
R6007 VSS.n2871 VSS.n2870 0.0147651
R6008 VSS.n3043 VSS.n2873 0.0147651
R6009 VSS.n1424 VSS.n1334 0.0147581
R6010 VSS.n1292 VSS.n9 0.0142813
R6011 VSS.n2929 VSS.n169 0.0140692
R6012 VSS.n2931 VSS.n177 0.0135154
R6013 VSS.n3007 VSS.n173 0.0135154
R6014 VSS.n3115 VSS.n3114 0.0124077
R6015 VSS.n3048 VSS.n168 0.0124077
R6016 VSS.n2854 VSS.t106 0.0121715
R6017 VSS.t107 VSS.n2874 0.0121715
R6018 VSS.n2952 VSS.n176 0.0118538
R6019 VSS.n972 VSS.n971 0.0115959
R6020 VSS.n3004 VSS.n173 0.0113
R6021 VSS.n3243 VSS.n119 0.0111996
R6022 VSS.n2841 VSS.n2836 0.011134
R6023 VSS.n3042 VSS.n2877 0.011134
R6024 VSS.n3426 VSS.n1 0.0110691
R6025 VSS.n3427 VSS.n3426 0.0110691
R6026 VSS.n3257 VSS.n107 0.0109186
R6027 VSS.n3094 VSS.n180 0.0107462
R6028 VSS.n3063 VSS.n167 0.0107462
R6029 VSS.n983 VSS.n982 0.0106712
R6030 VSS.n2970 VSS.n175 0.0101923
R6031 VSS.n976 VSS.n975 0.0100548
R6032 VSS.n957 VSS.n956 0.0100548
R6033 VSS.n3010 VSS.n3009 0.00978125
R6034 VSS.n3006 VSS.n2891 0.00978125
R6035 VSS.n2980 VSS.n174 0.00963846
R6036 VSS.n1417 VSS.n1382 0.00959535
R6037 VSS.n1465 VSS.n1454 0.00959535
R6038 VSS.n3082 VSS.n179 0.00908462
R6039 VSS.n2850 VSS.n179 0.00908462
R6040 VSS.n3044 VSS.t152 0.00854035
R6041 VSS.t152 VSS.n2869 0.00854035
R6042 VSS.n2989 VSS.n174 0.00853077
R6043 VSS.n3226 VSS.n3225 0.00833133
R6044 VSS.n3225 VSS.n3224 0.00833133
R6045 VSS.n3006 VSS.n105 0.00821305
R6046 VSS.n2967 VSS.n175 0.00797692
R6047 VSS.n3194 VSS.n109 0.00797126
R6048 VSS.t201 VSS.n109 0.00797126
R6049 VSS.n1117 VSS.n1114 0.00782743
R6050 VSS.n1419 VSS.n1418 0.00750352
R6051 VSS.n2830 VSS.n180 0.00742308
R6052 VSS.n3060 VSS.n167 0.00742308
R6053 VSS.n2841 VSS.t209 0.00655042
R6054 VSS.t106 VSS.n2841 0.00655042
R6055 VSS.n2871 VSS.t106 0.00655042
R6056 VSS.t152 VSS.n2871 0.00655042
R6057 VSS.t152 VSS.n3043 0.00655042
R6058 VSS.n3043 VSS.t107 0.00655042
R6059 VSS.t107 VSS.n3042 0.00655042
R6060 VSS.n3042 VSS.t108 0.00655042
R6061 VSS.n1373 VSS.n1372 0.00651467
R6062 VSS.n1371 VSS.n1297 0.00651467
R6063 VSS.n2942 VSS.n176 0.00631538
R6064 VSS.n3089 VSS.n2841 0.00594669
R6065 VSS.n3042 VSS.n2876 0.00594669
R6066 VSS.n3115 VSS.n181 0.00576154
R6067 VSS.n2919 VSS.n168 0.00576154
R6068 VSS.n1388 VSS.n1268 0.00554309
R6069 VSS.n1417 VSS.n1387 0.00554309
R6070 VSS.n1400 VSS.n1356 0.00554309
R6071 VSS.n1389 VSS.n1381 0.00554309
R6072 VSS.n1401 VSS.n1357 0.00554309
R6073 VSS.n1390 VSS.n1380 0.00554309
R6074 VSS.n1402 VSS.n1358 0.00554309
R6075 VSS.n1391 VSS.n1379 0.00554309
R6076 VSS.n1403 VSS.n1359 0.00554309
R6077 VSS.n1392 VSS.n1378 0.00554309
R6078 VSS.n1404 VSS.n1360 0.00554309
R6079 VSS.n1393 VSS.n1377 0.00554309
R6080 VSS.n1405 VSS.n1361 0.00554309
R6081 VSS.n1394 VSS.n1376 0.00554309
R6082 VSS.n1406 VSS.n1362 0.00554309
R6083 VSS.n1395 VSS.n1375 0.00554309
R6084 VSS.n1407 VSS.n1363 0.00554309
R6085 VSS.n1396 VSS.n1286 0.00554309
R6086 VSS.n1385 VSS.n1291 0.00554309
R6087 VSS.n1407 VSS.n1286 0.00554309
R6088 VSS.n1395 VSS.n1363 0.00554309
R6089 VSS.n1406 VSS.n1375 0.00554309
R6090 VSS.n1394 VSS.n1362 0.00554309
R6091 VSS.n1405 VSS.n1376 0.00554309
R6092 VSS.n1393 VSS.n1361 0.00554309
R6093 VSS.n1404 VSS.n1377 0.00554309
R6094 VSS.n1392 VSS.n1360 0.00554309
R6095 VSS.n1403 VSS.n1378 0.00554309
R6096 VSS.n1391 VSS.n1359 0.00554309
R6097 VSS.n1402 VSS.n1379 0.00554309
R6098 VSS.n1390 VSS.n1358 0.00554309
R6099 VSS.n1401 VSS.n1380 0.00554309
R6100 VSS.n1389 VSS.n1357 0.00554309
R6101 VSS.n1400 VSS.n1381 0.00554309
R6102 VSS.n1387 VSS.n1356 0.00554309
R6103 VSS.n1388 VSS.n1382 0.00554309
R6104 VSS.n1396 VSS.n1291 0.00554309
R6105 VSS.n1385 VSS.n1374 0.00554309
R6106 VSS.n1265 VSS.n1247 0.00554309
R6107 VSS.n1281 VSS.n1264 0.00554309
R6108 VSS.n1455 VSS.n1248 0.00554309
R6109 VSS.n1280 VSS.n1263 0.00554309
R6110 VSS.n1456 VSS.n1249 0.00554309
R6111 VSS.n1279 VSS.n1262 0.00554309
R6112 VSS.n1457 VSS.n1250 0.00554309
R6113 VSS.n1278 VSS.n1261 0.00554309
R6114 VSS.n1458 VSS.n1251 0.00554309
R6115 VSS.n1277 VSS.n1260 0.00554309
R6116 VSS.n1459 VSS.n1252 0.00554309
R6117 VSS.n1276 VSS.n1259 0.00554309
R6118 VSS.n1460 VSS.n1253 0.00554309
R6119 VSS.n1275 VSS.n1258 0.00554309
R6120 VSS.n1461 VSS.n1254 0.00554309
R6121 VSS.n1274 VSS.n1257 0.00554309
R6122 VSS.n1462 VSS.n1255 0.00554309
R6123 VSS.n1465 VSS.n1283 0.00554309
R6124 VSS.n1295 VSS.n1287 0.00554309
R6125 VSS.n1454 VSS.n1287 0.00554309
R6126 VSS.n1283 VSS.n1255 0.00554309
R6127 VSS.n1462 VSS.n1257 0.00554309
R6128 VSS.n1274 VSS.n1254 0.00554309
R6129 VSS.n1461 VSS.n1258 0.00554309
R6130 VSS.n1275 VSS.n1253 0.00554309
R6131 VSS.n1460 VSS.n1259 0.00554309
R6132 VSS.n1276 VSS.n1252 0.00554309
R6133 VSS.n1459 VSS.n1260 0.00554309
R6134 VSS.n1277 VSS.n1251 0.00554309
R6135 VSS.n1458 VSS.n1261 0.00554309
R6136 VSS.n1278 VSS.n1250 0.00554309
R6137 VSS.n1457 VSS.n1262 0.00554309
R6138 VSS.n1279 VSS.n1249 0.00554309
R6139 VSS.n1456 VSS.n1263 0.00554309
R6140 VSS.n1280 VSS.n1248 0.00554309
R6141 VSS.n1455 VSS.n1264 0.00554309
R6142 VSS.n1281 VSS.n1247 0.00554309
R6143 VSS.n1467 VSS.n1265 0.00554309
R6144 VSS.n1717 VSS.n1716 0.00508015
R6145 VSS.n1464 VSS.n1463 0.00507377
R6146 VSS.n1466 VSS.n1282 0.00507377
R6147 VSS.n3077 VSS.t106 0.00490922
R6148 VSS.t107 VSS.n2875 0.00490922
R6149 VSS VSS.n0 0.00466623
R6150 VSS.n2926 VSS.n177 0.00465385
R6151 VSS.n1082 VSS.n1076 0.0041
R6152 VSS.n2940 VSS.n169 0.0041
R6153 VSS.n1732 VSS.n1731 0.00405263
R6154 VSS.n901 VSS.n896 0.00405263
R6155 VSS.n1222 VSS.n1221 0.00372171
R6156 VSS.n1374 VSS.n1373 0.00358068
R6157 VSS.n1297 VSS.n1295 0.00358068
R6158 VSS.n3257 VSS.n3256 0.00338889
R6159 VSS.n3256 VSS.n3255 0.00338889
R6160 VSS.n1267 VSS.n1256 0.00328572
R6161 VSS.n1269 VSS.n1267 0.00328572
R6162 VSS.n1285 VSS.n1266 0.00328572
R6163 VSS.n1271 VSS.n1266 0.00328572
R6164 VSS.n1463 VSS.n1284 0.00328572
R6165 VSS.n1464 VSS.n1273 0.00328572
R6166 VSS.n1468 VSS.n1256 0.00328572
R6167 VSS.n1285 VSS.n1270 0.00328572
R6168 VSS.n1284 VSS.n1272 0.00328572
R6169 VSS.n1270 VSS.n1269 0.00328572
R6170 VSS.n1272 VSS.n1271 0.00328572
R6171 VSS.n1282 VSS.n1273 0.00328572
R6172 VSS.n949 VSS.n948 0.00327397
R6173 VSS.n3104 VSS.n165 0.00299231
R6174 VSS.n2859 VSS.n178 0.00299231
R6175 VSS.n1695 VSS.n1694 0.00296575
R6176 VSS.n1408 VSS.n1398 0.00296393
R6177 VSS.n1399 VSS.n1386 0.00296393
R6178 VSS.n1411 VSS.n1409 0.00296393
R6179 VSS.n1410 VSS.n1384 0.00296393
R6180 VSS.n1414 VSS.n1412 0.00296393
R6181 VSS.n1413 VSS.n1383 0.00296393
R6182 VSS.n1416 VSS.n1415 0.00296393
R6183 VSS.n1418 VSS.n1355 0.00296393
R6184 VSS.n1409 VSS.n1386 0.00296393
R6185 VSS.n1412 VSS.n1384 0.00296393
R6186 VSS.n1415 VSS.n1383 0.00296393
R6187 VSS.n1408 VSS.n1399 0.00296393
R6188 VSS.n1411 VSS.n1410 0.00296393
R6189 VSS.n1414 VSS.n1413 0.00296393
R6190 VSS.n1416 VSS.n1355 0.00296393
R6191 VSS.n1398 VSS.n1397 0.00296393
R6192 VSS.n3430 VSS.n1 0.00272514
R6193 VSS.n2906 VSS.n170 0.00243846
R6194 VSS.n2871 VSS.n2863 0.00231556
R6195 VSS.n3043 VSS.n2872 0.00231556
R6196 VSS.n3423 VSS.n1 0.00220437
R6197 VSS.n2991 VSS.n172 0.00188462
R6198 VSS.n2845 VSS.n166 0.00133077
R6199 VSS.n3109 VSS.t209 0.0012781
R6200 VSS.t108 VSS.n2880 0.0012781
R6201 VSS.n1712 VSS.n1711 0.00106849
R6202 VSS.t43 VSS.n1419 0.00100704
R6203 VSS.n2978 VSS.n171 0.000776923
R6204 VSS.n1118 VSS.n1072 0.000659292
R6205 VDD.n414 VDD.t265 589.355
R6206 VDD.n413 VDD.t218 589.355
R6207 VDD.n407 VDD.t231 589.355
R6208 VDD.n400 VDD.t227 589.355
R6209 VDD.n393 VDD.t222 589.355
R6210 VDD.n386 VDD.t237 589.355
R6211 VDD.n379 VDD.t220 589.355
R6212 VDD.n372 VDD.t229 589.355
R6213 VDD.n208 VDD.t306 484.969
R6214 VDD.t302 VDD.n207 480.769
R6215 VDD.n186 VDD.t102 448.111
R6216 VDD.n198 VDD.t253 443.911
R6217 VDD.t282 VDD.n198 443.911
R6218 VDD.n199 VDD.t35 443.911
R6219 VDD.n199 VDD.t280 443.911
R6220 VDD.n207 VDD.t280 443.911
R6221 VDD.n408 VDD.t189 419.211
R6222 VDD.n401 VDD.t95 419.211
R6223 VDD.n394 VDD.t41 419.211
R6224 VDD.n387 VDD.t249 419.211
R6225 VDD.n380 VDD.t28 419.211
R6226 VDD.n373 VDD.t215 419.211
R6227 VDD.t19 VDD.t82 416.988
R6228 VDD.t224 VDD.t267 403.476
R6229 VDD.t25 VDD.t2 384.764
R6230 VDD.t16 VDD.t47 372.587
R6231 VDD.t247 VDD.t39 372.228
R6232 VDD.t23 VDD.t91 372.228
R6233 VDD.t304 VDD.t302 346.154
R6234 VDD.t107 VDD.t304 346.154
R6235 VDD.t306 VDD.t107 346.154
R6236 VDD.n127 VDD.t33 345.56
R6237 VDD.t33 VDD.t132 335.908
R6238 VDD.n128 VDD.t134 320.464
R6239 VDD.t88 VDD.t4 288.611
R6240 VDD.t286 VDD.t98 282.546
R6241 VDD.n117 VDD.t187 282.116
R6242 VDD.n141 VDD.t49 282.116
R6243 VDD.n83 VDD.t139 281.861
R6244 VDD.t114 VDD.n147 279.923
R6245 VDD.n146 VDD.t12 278.959
R6246 VDD.t272 VDD.t96 277.027
R6247 VDD.t18 VDD.t88 275.098
R6248 VDD.t102 VDD.t308 272.437
R6249 VDD.t308 VDD.t37 272.437
R6250 VDD.t37 VDD.t284 272.437
R6251 VDD.t284 VDD.t15 272.437
R6252 VDD.t15 VDD.t106 272.437
R6253 VDD.t106 VDD.t14 272.437
R6254 VDD.t14 VDD.t44 272.437
R6255 VDD.t44 VDD.t260 272.437
R6256 VDD.t260 VDD.t259 272.437
R6257 VDD.t259 VDD.t257 272.437
R6258 VDD.t257 VDD.t258 272.437
R6259 VDD.t258 VDD.t136 272.437
R6260 VDD.t136 VDD.t300 272.437
R6261 VDD.t300 VDD.t42 272.437
R6262 VDD.t42 VDD.t253 272.437
R6263 VDD.t137 VDD.t282 272.437
R6264 VDD.t285 VDD.t137 272.437
R6265 VDD.t35 VDD.t285 272.437
R6266 VDD.t132 VDD.t31 239.382
R6267 VDD.t113 VDD.t10 238.188
R6268 VDD.t66 VDD.t76 235.522
R6269 VDD.t183 VDD.t199 235.522
R6270 VDD.n95 VDD.t80 233.591
R6271 VDD.t68 VDD.t235 231.661
R6272 VDD.t261 VDD.n145 224.436
R6273 VDD.n81 VDD.t164 219.865
R6274 VDD.n151 VDD.n150 217.452
R6275 VDD.t151 VDD.t155 216.216
R6276 VDD.t29 VDD.n81 212.15
R6277 VDD.t298 VDD.t173 211.391
R6278 VDD.t4 VDD.t0 208.494
R6279 VDD.n34 VDD.n6 199.776
R6280 VDD.n34 VDD.n7 199.776
R6281 VDD.n32 VDD.n6 199.776
R6282 VDD.n32 VDD.n7 199.776
R6283 VDD.n46 VDD.n40 199.776
R6284 VDD.n46 VDD.n41 199.776
R6285 VDD.n44 VDD.n40 199.776
R6286 VDD.n44 VDD.n41 199.776
R6287 VDD.t8 VDD.t276 196.911
R6288 VDD.t89 VDD.t274 196.911
R6289 VDD.t274 VDD.t62 196.911
R6290 VDD.t111 VDD.t60 196.911
R6291 VDD.t244 VDD.t290 196.911
R6292 VDD.t82 VDD.t224 196.911
R6293 VDD.t70 VDD.t74 196.911
R6294 VDD.t292 VDD.t255 196.721
R6295 VDD.t296 VDD.t6 196.721
R6296 VDD.t93 VDD.t126 196.721
R6297 VDD.n34 VDD.t239 187.815
R6298 VDD.t216 VDD.n32 187.815
R6299 VDD.n46 VDD.t193 187.815
R6300 VDD.t157 VDD.n44 187.815
R6301 VDD.t251 VDD.t153 181.468
R6302 VDD.t21 VDD.t244 174.71
R6303 VDD.t126 VDD.t318 174.542
R6304 VDD.t169 VDD.t72 173.745
R6305 VDD.t60 VDD.t21 168.919
R6306 VDD.t318 VDD.t296 168.756
R6307 VDD.t58 VDD.t84 167.954
R6308 VDD.t199 VDD.t116 167.954
R6309 VDD.t204 VDD.t151 166.024
R6310 VDD.t294 VDD.t64 162.162
R6311 VDD.n60 VDD.t288 156.802
R6312 VDD.t45 VDD.t272 155.405
R6313 VDD.n147 VDD.t58 152.511
R6314 VDD.t31 VDD.t18 150.579
R6315 VDD.t53 VDD.t203 150.579
R6316 VDD.t104 VDD.t292 149.47
R6317 VDD.t181 VDD.t286 149.47
R6318 VDD.t0 VDD.t86 142.857
R6319 VDD.t51 VDD.t138 142.857
R6320 VDD.n126 VDD.t19 138.031
R6321 VDD.t74 VDD.t100 121.623
R6322 VDD.t80 VDD.t55 119.692
R6323 VDD.t130 VDD.t233 119.692
R6324 VDD.t100 VDD.t78 113.9
R6325 VDD.t84 VDD.n146 111.969
R6326 VDD.t239 VDD.t176 107.053
R6327 VDD.t176 VDD.t243 107.053
R6328 VDD.t243 VDD.t212 107.053
R6329 VDD.t212 VDD.t179 107.053
R6330 VDD.t179 VDD.t178 107.053
R6331 VDD.t178 VDD.t217 107.053
R6332 VDD.t217 VDD.t269 107.053
R6333 VDD.t269 VDD.t177 107.053
R6334 VDD.t177 VDD.t315 107.053
R6335 VDD.t214 VDD.t213 107.053
R6336 VDD.t213 VDD.t180 107.053
R6337 VDD.t180 VDD.t240 107.053
R6338 VDD.t240 VDD.t271 107.053
R6339 VDD.t271 VDD.t270 107.053
R6340 VDD.t270 VDD.t316 107.053
R6341 VDD.t316 VDD.t242 107.053
R6342 VDD.t242 VDD.t241 107.053
R6343 VDD.t241 VDD.t216 107.053
R6344 VDD.t193 VDD.t194 107.053
R6345 VDD.t194 VDD.t299 107.053
R6346 VDD.t299 VDD.t142 107.053
R6347 VDD.t142 VDD.t313 107.053
R6348 VDD.t313 VDD.t163 107.053
R6349 VDD.t163 VDD.t202 107.053
R6350 VDD.t202 VDD.t195 107.053
R6351 VDD.t195 VDD.t158 107.053
R6352 VDD.t158 VDD.t160 107.053
R6353 VDD.t175 VDD.t312 107.053
R6354 VDD.t312 VDD.t196 107.053
R6355 VDD.t196 VDD.t161 107.053
R6356 VDD.t161 VDD.t141 107.053
R6357 VDD.t141 VDD.t166 107.053
R6358 VDD.t166 VDD.t162 107.053
R6359 VDD.t162 VDD.t201 107.053
R6360 VDD.t201 VDD.t159 107.053
R6361 VDD.t159 VDD.t157 107.053
R6362 VDD.t288 VDD.t113 98.3612
R6363 VDD.t233 VDD.t51 88.8036
R6364 VDD.n94 VDD.t149 87.8383
R6365 VDD.t255 VDD.t247 85.825
R6366 VDD.t55 VDD.t66 77.2206
R6367 VDD.t173 VDD.t130 77.2206
R6368 VDD.t86 VDD.n126 71.4291
R6369 VDD.t171 VDD.n94 67.5681
R6370 VDD.n245 VDD.n244 66.6672
R6371 VDD.n257 VDD.n231 66.6672
R6372 VDD.n259 VDD.n258 66.6672
R6373 VDD.n271 VDD.n223 66.6672
R6374 VDD.n273 VDD.n272 66.6672
R6375 VDD.n286 VDD.n215 66.6672
R6376 VDD.n288 VDD.n287 66.6672
R6377 VDD.t96 VDD.t111 66.6028
R6378 VDD.n361 VDD.n360 66.5439
R6379 VDD.n359 VDD.n314 66.5439
R6380 VDD.n351 VDD.n350 66.5439
R6381 VDD.n349 VDD.n318 66.5439
R6382 VDD.n341 VDD.n340 66.5439
R6383 VDD.n339 VDD.n322 66.5439
R6384 VDD.n331 VDD.n330 66.5439
R6385 VDD.t6 VDD.t29 66.5386
R6386 VDD.t128 VDD.n243 66.177
R6387 VDD.t143 VDD.n311 66.0664
R6388 VDD.t72 VDD.t53 65.6376
R6389 VDD.n17 VDD.n15 65.4873
R6390 VDD.n20 VDD.n14 65.4873
R6391 VDD.t290 VDD.t16 60.8113
R6392 VDD.t98 VDD.t93 60.7527
R6393 VDD.n245 VDD.t124 59.877
R6394 VDD.t190 VDD.n257 59.877
R6395 VDD.n259 VDD.t118 59.877
R6396 VDD.t185 VDD.n271 59.877
R6397 VDD.n273 VDD.t120 59.877
R6398 VDD.t310 VDD.n286 59.877
R6399 VDD.n288 VDD.t122 59.877
R6400 VDD.t47 VDD.t261 59.8461
R6401 VDD.t39 VDD.t23 59.7883
R6402 VDD.t91 VDD.t164 59.7883
R6403 VDD.n360 VDD.t208 59.7664
R6404 VDD.t147 VDD.n314 59.7664
R6405 VDD.n350 VDD.t197 59.7664
R6406 VDD.t145 VDD.n318 59.7664
R6407 VDD.n340 VDD.t109 59.7664
R6408 VDD.t206 VDD.n322 59.7664
R6409 VDD.n330 VDD.t210 59.7664
R6410 VDD.n150 VDD.t8 56.9503
R6411 VDD.t315 VDD.n33 53.527
R6412 VDD.n33 VDD.t214 53.527
R6413 VDD.t160 VDD.n45 53.527
R6414 VDD.n45 VDD.t175 53.527
R6415 VDD.t149 VDD.t204 50.1936
R6416 VDD.t267 VDD.t49 48.263
R6417 VDD.t116 VDD.t187 48.263
R6418 VDD.t139 VDD.t25 48.2165
R6419 VDD.n18 VDD.n14 48.0418
R6420 VDD.n19 VDD.n15 48.0418
R6421 VDD.t10 VDD.t104 47.2522
R6422 VDD.t2 VDD.t181 47.2522
R6423 VDD.n151 VDD.t278 44.4358
R6424 VDD.t12 VDD.t45 41.5063
R6425 VDD.t276 VDD.t294 34.7495
R6426 VDD.t64 VDD.t89 34.7495
R6427 VDD.t155 VDD.t251 34.7495
R6428 VDD.t62 VDD.t114 29.9233
R6429 VDD.t235 VDD.t298 24.1318
R6430 VDD.t76 VDD.t169 23.1665
R6431 VDD.n135 VDD.t57 21.6375
R6432 VDD.n135 VDD.t20 21.6375
R6433 VDD.n109 VDD.t205 21.6375
R6434 VDD.t203 VDD.t68 19.3055
R6435 VDD.n94 VDD.t27 16.2012
R6436 VDD.n126 VDD.t246 15.981
R6437 VDD.t153 VDD.t183 15.4445
R6438 VDD.n201 VDD.t281 12.2195
R6439 VDD.n291 VDD.t122 12.1776
R6440 VDD.t210 VDD.n329 12.1637
R6441 VDD.n292 VDD.n291 11.4951
R6442 VDD.n329 VDD.n326 11.4938
R6443 VDD.n207 VDD.n206 11.0111
R6444 VDD.n200 VDD.n199 11.0111
R6445 VDD.n198 VDD.n197 11.0111
R6446 VDD.n185 VDD.t36 10.0145
R6447 VDD.n196 VDD.t283 10.0145
R6448 VDD.n195 VDD.t254 10.0145
R6449 VDD.n202 VDD.t307 9.42355
R6450 VDD.n205 VDD.t303 9.42355
R6451 VDD.n194 VDD.n193 8.54446
R6452 VDD.n192 VDD.n191 8.54446
R6453 VDD.n414 VDD.t266 8.52192
R6454 VDD.n413 VDD.t219 8.52192
R6455 VDD.n407 VDD.t232 8.46717
R6456 VDD.n400 VDD.t228 8.46717
R6457 VDD.n393 VDD.t223 8.46717
R6458 VDD.n386 VDD.t238 8.46717
R6459 VDD.n379 VDD.t221 8.46717
R6460 VDD.n372 VDD.t230 8.46717
R6461 VDD.n204 VDD.n203 8.11105
R6462 VDD.n128 VDD.n127 7.72251
R6463 VDD VDD.n417 7.7195
R6464 VDD.n115 VDD.t188 7.51784
R6465 VDD.n107 VDD.t172 7.5061
R6466 VDD.n155 VDD.t295 7.46
R6467 VDD.n158 VDD.t63 7.46
R6468 VDD.n125 VDD.t264 7.40883
R6469 VDD.n124 VDD.t32 7.40883
R6470 VDD.n91 VDD.t54 7.40883
R6471 VDD.n244 VDD.t128 6.79062
R6472 VDD.t124 VDD.n231 6.79062
R6473 VDD.n258 VDD.t190 6.79062
R6474 VDD.t118 VDD.n223 6.79062
R6475 VDD.n272 VDD.t185 6.79062
R6476 VDD.t120 VDD.n215 6.79062
R6477 VDD.n287 VDD.t310 6.79062
R6478 VDD.n361 VDD.t143 6.77807
R6479 VDD.t208 VDD.n359 6.77807
R6480 VDD.n351 VDD.t147 6.77807
R6481 VDD.t197 VDD.n349 6.77807
R6482 VDD.n341 VDD.t145 6.77807
R6483 VDD.t109 VDD.n339 6.77807
R6484 VDD.n331 VDD.t206 6.77807
R6485 VDD.n290 VDD.n211 6.3005
R6486 VDD.n289 VDD.n214 6.3005
R6487 VDD.n289 VDD.n288 6.3005
R6488 VDD.n219 VDD.n212 6.3005
R6489 VDD.n287 VDD.n212 6.3005
R6490 VDD.n285 VDD.n284 6.3005
R6491 VDD.n286 VDD.n285 6.3005
R6492 VDD.n277 VDD.n216 6.3005
R6493 VDD.n216 VDD.n215 6.3005
R6494 VDD.n275 VDD.n274 6.3005
R6495 VDD.n274 VDD.n273 6.3005
R6496 VDD.n227 VDD.n222 6.3005
R6497 VDD.n272 VDD.n222 6.3005
R6498 VDD.n270 VDD.n269 6.3005
R6499 VDD.n271 VDD.n270 6.3005
R6500 VDD.n263 VDD.n224 6.3005
R6501 VDD.n224 VDD.n223 6.3005
R6502 VDD.n261 VDD.n260 6.3005
R6503 VDD.n260 VDD.n259 6.3005
R6504 VDD.n235 VDD.n230 6.3005
R6505 VDD.n258 VDD.n230 6.3005
R6506 VDD.n256 VDD.n255 6.3005
R6507 VDD.n257 VDD.n256 6.3005
R6508 VDD.n249 VDD.n232 6.3005
R6509 VDD.n232 VDD.n231 6.3005
R6510 VDD.n247 VDD.n246 6.3005
R6511 VDD.n246 VDD.n245 6.3005
R6512 VDD.n239 VDD.n238 6.3005
R6513 VDD.n244 VDD.n238 6.3005
R6514 VDD.n243 VDD.n242 6.3005
R6515 VDD.n311 VDD.n310 6.3005
R6516 VDD.n363 VDD.n362 6.3005
R6517 VDD.n362 VDD.n361 6.3005
R6518 VDD.n313 VDD.n312 6.3005
R6519 VDD.n360 VDD.n313 6.3005
R6520 VDD.n358 VDD.n357 6.3005
R6521 VDD.n359 VDD.n358 6.3005
R6522 VDD.n356 VDD.n355 6.3005
R6523 VDD.n356 VDD.n314 6.3005
R6524 VDD.n352 VDD.n317 6.3005
R6525 VDD.n352 VDD.n351 6.3005
R6526 VDD.n316 VDD.n315 6.3005
R6527 VDD.n350 VDD.n316 6.3005
R6528 VDD.n348 VDD.n347 6.3005
R6529 VDD.n349 VDD.n348 6.3005
R6530 VDD.n346 VDD.n345 6.3005
R6531 VDD.n346 VDD.n318 6.3005
R6532 VDD.n342 VDD.n321 6.3005
R6533 VDD.n342 VDD.n341 6.3005
R6534 VDD.n320 VDD.n319 6.3005
R6535 VDD.n340 VDD.n320 6.3005
R6536 VDD.n338 VDD.n337 6.3005
R6537 VDD.n339 VDD.n338 6.3005
R6538 VDD.n336 VDD.n335 6.3005
R6539 VDD.n336 VDD.n322 6.3005
R6540 VDD.n332 VDD.n325 6.3005
R6541 VDD.n332 VDD.n331 6.3005
R6542 VDD.n324 VDD.n323 6.3005
R6543 VDD.n330 VDD.n324 6.3005
R6544 VDD.n328 VDD.n327 6.3005
R6545 VDD.n123 VDD.t317 6.22272
R6546 VDD.n122 VDD.t1 6.22272
R6547 VDD.n88 VDD.t52 6.22272
R6548 VDD.n417 VDD.n416 6.1835
R6549 VDD.n417 VDD.n56 6.09991
R6550 VDD.n243 VDD.n238 6.0755
R6551 VDD.n246 VDD.n238 6.0755
R6552 VDD.n246 VDD.n232 6.0755
R6553 VDD.n256 VDD.n232 6.0755
R6554 VDD.n256 VDD.n230 6.0755
R6555 VDD.n260 VDD.n230 6.0755
R6556 VDD.n260 VDD.n224 6.0755
R6557 VDD.n270 VDD.n224 6.0755
R6558 VDD.n270 VDD.n222 6.0755
R6559 VDD.n274 VDD.n222 6.0755
R6560 VDD.n274 VDD.n216 6.0755
R6561 VDD.n285 VDD.n216 6.0755
R6562 VDD.n285 VDD.n212 6.0755
R6563 VDD.n289 VDD.n212 6.0755
R6564 VDD.n290 VDD.n289 6.0755
R6565 VDD.n362 VDD.n311 6.0755
R6566 VDD.n362 VDD.n313 6.0755
R6567 VDD.n358 VDD.n313 6.0755
R6568 VDD.n358 VDD.n356 6.0755
R6569 VDD.n356 VDD.n352 6.0755
R6570 VDD.n352 VDD.n316 6.0755
R6571 VDD.n348 VDD.n316 6.0755
R6572 VDD.n348 VDD.n346 6.0755
R6573 VDD.n346 VDD.n342 6.0755
R6574 VDD.n342 VDD.n320 6.0755
R6575 VDD.n338 VDD.n320 6.0755
R6576 VDD.n338 VDD.n336 6.0755
R6577 VDD.n336 VDD.n332 6.0755
R6578 VDD.n332 VDD.n324 6.0755
R6579 VDD.n328 VDD.n324 6.0755
R6580 VDD.n133 VDD.n124 5.49789
R6581 VDD.n133 VDD.n125 5.49789
R6582 VDD.n103 VDD.n91 5.49789
R6583 VDD.n134 VDD.n122 5.41359
R6584 VDD.n134 VDD.n123 5.41359
R6585 VDD.n106 VDD.n88 5.41359
R6586 VDD.n110 VDD.n87 5.35702
R6587 VDD.n105 VDD.n89 5.35702
R6588 VDD.n102 VDD.n92 5.35702
R6589 VDD.n100 VDD.n93 5.35702
R6590 VDD.n98 VDD.n96 5.35702
R6591 VDD.n136 VDD.n120 5.35271
R6592 VDD.n136 VDD.n121 5.35271
R6593 VDD.n111 VDD.n86 5.35271
R6594 VDD.n112 VDD.n85 5.31398
R6595 VDD.n157 VDD.n148 5.30615
R6596 VDD.n154 VDD.n149 5.29976
R6597 VDD.n62 VDD.n59 5.29976
R6598 VDD.n104 VDD.n90 5.28659
R6599 VDD.n123 VDD.t5 5.05606
R6600 VDD.n122 VDD.t250 5.05606
R6601 VDD.n88 VDD.t131 5.05606
R6602 VDD.n38 VDD.n37 4.94375
R6603 VDD VDD.n0 4.82228
R6604 VDD.n156 VDD.t65 4.70061
R6605 VDD.n64 VDD.t256 4.70061
R6606 VDD.n241 VDD.n240 4.60502
R6607 VDD.n209 VDD.n208 4.56013
R6608 VDD.n208 VDD.n57 4.56013
R6609 VDD.n202 VDD.n184 4.55193
R6610 VDD.n409 VDD.n406 4.5005
R6611 VDD.n406 VDD.n405 4.5005
R6612 VDD.n409 VDD.n408 4.5005
R6613 VDD.n408 VDD.n405 4.5005
R6614 VDD.n402 VDD.n399 4.5005
R6615 VDD.n399 VDD.n398 4.5005
R6616 VDD.n402 VDD.n401 4.5005
R6617 VDD.n401 VDD.n398 4.5005
R6618 VDD.n395 VDD.n392 4.5005
R6619 VDD.n392 VDD.n391 4.5005
R6620 VDD.n395 VDD.n394 4.5005
R6621 VDD.n394 VDD.n391 4.5005
R6622 VDD.n388 VDD.n385 4.5005
R6623 VDD.n385 VDD.n384 4.5005
R6624 VDD.n388 VDD.n387 4.5005
R6625 VDD.n387 VDD.n384 4.5005
R6626 VDD.n381 VDD.n378 4.5005
R6627 VDD.n378 VDD.n377 4.5005
R6628 VDD.n381 VDD.n380 4.5005
R6629 VDD.n380 VDD.n377 4.5005
R6630 VDD.n374 VDD.n371 4.5005
R6631 VDD.n371 VDD.n370 4.5005
R6632 VDD.n374 VDD.n373 4.5005
R6633 VDD.n373 VDD.n370 4.5005
R6634 VDD.n24 VDD.n23 4.5005
R6635 VDD.n30 VDD.n29 4.5005
R6636 VDD.n28 VDD.n10 4.5005
R6637 VDD.n27 VDD.n26 4.5005
R6638 VDD.n25 VDD.n11 4.5005
R6639 VDD.n53 VDD.n1 4.5005
R6640 VDD.n52 VDD.n51 4.5005
R6641 VDD.n50 VDD.n3 4.5005
R6642 VDD.n49 VDD.n48 4.5005
R6643 VDD.n55 VDD.n54 4.5005
R6644 VDD.n294 VDD.n293 4.5005
R6645 VDD.n213 VDD.n210 4.5005
R6646 VDD.n281 VDD.n280 4.5005
R6647 VDD.n283 VDD.n282 4.5005
R6648 VDD.n279 VDD.n278 4.5005
R6649 VDD.n276 VDD.n220 4.5005
R6650 VDD.n266 VDD.n221 4.5005
R6651 VDD.n268 VDD.n267 4.5005
R6652 VDD.n265 VDD.n264 4.5005
R6653 VDD.n262 VDD.n228 4.5005
R6654 VDD.n252 VDD.n229 4.5005
R6655 VDD.n254 VDD.n253 4.5005
R6656 VDD.n251 VDD.n250 4.5005
R6657 VDD.n248 VDD.n236 4.5005
R6658 VDD.n240 VDD.n237 4.5005
R6659 VDD.n182 VDD.n58 4.5005
R6660 VDD.n365 VDD.n302 4.5005
R6661 VDD.n365 VDD.n303 4.5005
R6662 VDD.n365 VDD.n301 4.5005
R6663 VDD.n365 VDD.n304 4.5005
R6664 VDD.n365 VDD.n300 4.5005
R6665 VDD.n365 VDD.n305 4.5005
R6666 VDD.n365 VDD.n299 4.5005
R6667 VDD.n365 VDD.n306 4.5005
R6668 VDD.n365 VDD.n298 4.5005
R6669 VDD.n365 VDD.n307 4.5005
R6670 VDD.n365 VDD.n297 4.5005
R6671 VDD.n365 VDD.n308 4.5005
R6672 VDD.n365 VDD.n296 4.5005
R6673 VDD.n365 VDD.n309 4.5005
R6674 VDD.n365 VDD.n295 4.5005
R6675 VDD.n365 VDD.n364 4.5005
R6676 VDD.n189 VDD.n186 4.5005
R6677 VDD.n189 VDD.n188 4.5005
R6678 VDD.n172 VDD.t291 4.46351
R6679 VDD.n170 VDD.t245 4.46351
R6680 VDD.n169 VDD.t61 4.46351
R6681 VDD.n167 VDD.t112 4.46351
R6682 VDD.n166 VDD.t273 4.46351
R6683 VDD.n164 VDD.t13 4.46351
R6684 VDD.n70 VDD.t3 4.46351
R6685 VDD.n72 VDD.t287 4.46351
R6686 VDD.n73 VDD.t94 4.46351
R6687 VDD.n75 VDD.t127 4.46351
R6688 VDD.n76 VDD.t297 4.46351
R6689 VDD.n78 VDD.t7 4.46351
R6690 VDD.n129 VDD.t192 4.45405
R6691 VDD.n97 VDD.t79 4.385
R6692 VDD.n175 VDD.t48 4.36426
R6693 VDD.n161 VDD.t59 4.36426
R6694 VDD.n159 VDD.t115 4.36426
R6695 VDD.n152 VDD.t279 4.36426
R6696 VDD.n139 VDD.t50 4.36426
R6697 VDD.n82 VDD.t140 4.36426
R6698 VDD.n68 VDD.t92 4.36426
R6699 VDD.n66 VDD.t40 4.36426
R6700 VDD.n60 VDD.t289 4.36426
R6701 VDD.n163 VDD.t85 4.36035
R6702 VDD.n165 VDD.t46 4.36035
R6703 VDD.n168 VDD.t97 4.36035
R6704 VDD.n171 VDD.t22 4.36035
R6705 VDD.n173 VDD.t17 4.36035
R6706 VDD.n177 VDD.t262 4.36035
R6707 VDD.n129 VDD.t135 4.36035
R6708 VDD.n137 VDD.t268 4.36035
R6709 VDD.n97 VDD.t101 4.36035
R6710 VDD.n113 VDD.t117 4.36035
R6711 VDD.n61 VDD.t105 4.36035
R6712 VDD.n63 VDD.t248 4.36035
R6713 VDD.n65 VDD.t24 4.36035
R6714 VDD.n67 VDD.t165 4.36035
R6715 VDD.n79 VDD.t30 4.36035
R6716 VDD.n77 VDD.t319 4.36035
R6717 VDD.n74 VDD.t99 4.36035
R6718 VDD.n71 VDD.t182 4.36035
R6719 VDD.n69 VDD.t26 4.36035
R6720 VDD.n162 VDD.n146 4.35926
R6721 VDD.n131 VDD.n127 4.35926
R6722 VDD.n81 VDD.n80 4.35926
R6723 VDD.n153 VDD.n150 4.35925
R6724 VDD.n160 VDD.n147 4.35925
R6725 VDD.n130 VDD.n128 4.35925
R6726 VDD.n99 VDD.n95 4.35925
R6727 VDD.n132 VDD.t263 4.29774
R6728 VDD.n132 VDD.t34 4.29774
R6729 VDD.n101 VDD.t56 4.29774
R6730 VDD.n108 VDD.t150 4.28209
R6731 VDD.n23 VDD.n22 4.1815
R6732 VDD.n85 VDD.t154 3.91054
R6733 VDD.t138 VDD.t171 3.8615
R6734 VDD.n90 VDD.t236 3.7566
R6735 VDD.n188 VDD.t103 3.20383
R6736 VDD.n152 VDD.n151 3.05229
R6737 VDD.n369 VDD.n182 2.97032
R6738 VDD.n43 VDD.n42 2.85445
R6739 VDD.n43 VDD.n2 2.85445
R6740 VDD.n369 VDD.n57 2.82015
R6741 VDD.n411 VDD.n410 2.70462
R6742 VDD.n404 VDD.n403 2.70462
R6743 VDD.n397 VDD.n396 2.70462
R6744 VDD.n390 VDD.n389 2.70462
R6745 VDD.n383 VDD.n382 2.70462
R6746 VDD.n376 VDD.n375 2.70462
R6747 VDD.n9 VDD.n8 2.5272
R6748 VDD.n8 VDD.n4 2.5272
R6749 VDD.n36 VDD.n5 2.5272
R6750 VDD.n42 VDD.n39 2.5272
R6751 VDD.n192 VDD.n190 2.38453
R6752 VDD.n179 VDD.n145 2.29149
R6753 VDD.n24 VDD.n5 2.28609
R6754 VDD.n54 VDD.n2 2.28609
R6755 VDD.n174 VDD.n144 2.28317
R6756 VDD.n138 VDD.n119 2.28317
R6757 VDD.n114 VDD.n84 2.28317
R6758 VDD.n125 VDD.t133 2.2755
R6759 VDD.n124 VDD.t314 2.2755
R6760 VDD.n91 VDD.t170 2.2755
R6761 VDD.n416 VDD.n415 2.25109
R6762 VDD.n179 VDD.n178 2.2505
R6763 VDD.n176 VDD.n144 2.2505
R6764 VDD.n140 VDD.n119 2.2505
R6765 VDD.n116 VDD.n84 2.2505
R6766 VDD.n187 VDD.n0 2.23822
R6767 VDD.n85 VDD.t200 2.22001
R6768 VDD.n89 VDD.t174 2.22001
R6769 VDD.n89 VDD.t234 2.22001
R6770 VDD.n148 VDD.t90 2.15435
R6771 VDD.n148 VDD.t275 2.15435
R6772 VDD.n121 VDD.t87 2.10455
R6773 VDD.n121 VDD.t225 2.10455
R6774 VDD.n120 VDD.t83 2.10455
R6775 VDD.n120 VDD.t226 2.10455
R6776 VDD.n86 VDD.t252 2.10455
R6777 VDD.n86 VDD.t184 2.10455
R6778 VDD.n87 VDD.t152 2.06607
R6779 VDD.n310 VDD.t144 2.04514
R6780 VDD.n242 VDD.t129 2.04159
R6781 VDD.n56 VDD.n55 2.02679
R6782 VDD.n326 VDD.t211 2.02385
R6783 VDD.n13 VDD.t168 2.0205
R6784 VDD.n292 VDD.t123 2.0203
R6785 VDD.n95 VDD.t70 1.931
R6786 VDD.n412 VDD.n56 1.88697
R6787 VDD.n149 VDD.t9 1.84822
R6788 VDD.n149 VDD.t277 1.84822
R6789 VDD.n59 VDD.t11 1.84822
R6790 VDD.n59 VDD.t293 1.84822
R6791 VDD.n416 VDD.n412 1.81813
R6792 VDD.n90 VDD.t69 1.67844
R6793 VDD.n21 VDD.n20 1.5755
R6794 VDD.n17 VDD.n16 1.5755
R6795 VDD.n87 VDD.t156 1.4923
R6796 VDD.n92 VDD.t77 1.4923
R6797 VDD.n92 VDD.t73 1.4923
R6798 VDD.n93 VDD.t81 1.4923
R6799 VDD.n93 VDD.t67 1.4923
R6800 VDD.n96 VDD.t75 1.4923
R6801 VDD.n96 VDD.t71 1.4923
R6802 VDD.n182 VDD.n83 1.48949
R6803 VDD.n334 VDD.n333 1.47853
R6804 VDD.n344 VDD.n343 1.47853
R6805 VDD.n354 VDD.n353 1.47853
R6806 VDD.n234 VDD.n233 1.47497
R6807 VDD.n226 VDD.n225 1.47497
R6808 VDD.n218 VDD.n217 1.47497
R6809 VDD.n182 VDD.n181 1.46788
R6810 VDD.n383 VDD.n376 1.4375
R6811 VDD.n390 VDD.n383 1.4375
R6812 VDD.n397 VDD.n390 1.4375
R6813 VDD.n404 VDD.n397 1.4375
R6814 VDD.n411 VDD.n404 1.4375
R6815 VDD.n412 VDD.n411 1.4375
R6816 VDD.n19 VDD.t167 1.15641
R6817 VDD.t167 VDD.n18 1.15641
R6818 VDD.n142 VDD.n141 1.14644
R6819 VDD.n118 VDD.n117 1.14644
R6820 VDD.n29 VDD.n9 1.06648
R6821 VDD.n366 VDD.n183 1.02433
R6822 VDD.n37 VDD.n4 1.00685
R6823 VDD.n37 VDD.n36 1.00685
R6824 VDD.n39 VDD.n38 1.00685
R6825 VDD.n16 VDD.n12 0.936026
R6826 VDD.n143 VDD.n118 0.9215
R6827 VDD.n193 VDD.t301 0.9105
R6828 VDD.n193 VDD.t43 0.9105
R6829 VDD.n191 VDD.t309 0.9105
R6830 VDD.n191 VDD.t38 0.9105
R6831 VDD.n203 VDD.t305 0.813
R6832 VDD.n203 VDD.t108 0.813
R6833 VDD.n14 VDD.n13 0.788
R6834 VDD.n15 VDD.n12 0.788
R6835 VDD.n32 VDD.n31 0.788
R6836 VDD.n35 VDD.n34 0.788
R6837 VDD.n44 VDD.n43 0.788
R6838 VDD.n47 VDD.n46 0.788
R6839 VDD.n367 VDD.n294 0.7505
R6840 VDD.n21 VDD.n13 0.734526
R6841 VDD.n16 VDD.n13 0.734526
R6842 VDD.n22 VDD.n12 0.676711
R6843 VDD.n194 VDD.n192 0.656214
R6844 VDD.n143 VDD.n142 0.563
R6845 VDD.n181 VDD.n180 0.563
R6846 VDD.n368 VDD.n183 0.555536
R6847 VDD.n367 VDD.n366 0.54104
R6848 VDD.n329 VDD.n328 0.450111
R6849 VDD.n291 VDD.n290 0.449462
R6850 VDD.n18 VDD.n17 0.410734
R6851 VDD.n20 VDD.n19 0.410734
R6852 VDD.n376 VDD.n369 0.386525
R6853 VDD.n181 VDD.n143 0.359
R6854 VDD.n233 VDD.t125 0.3255
R6855 VDD.n233 VDD.t191 0.3255
R6856 VDD.n225 VDD.t119 0.3255
R6857 VDD.n225 VDD.t186 0.3255
R6858 VDD.n217 VDD.t121 0.3255
R6859 VDD.n217 VDD.t311 0.3255
R6860 VDD.n333 VDD.t110 0.3255
R6861 VDD.n333 VDD.t207 0.3255
R6862 VDD.n343 VDD.t198 0.3255
R6863 VDD.n343 VDD.t146 0.3255
R6864 VDD.n353 VDD.t209 0.3255
R6865 VDD.n353 VDD.t148 0.3255
R6866 VDD.n134 VDD.n133 0.305021
R6867 VDD.n31 VDD.n9 0.272055
R6868 VDD.n35 VDD.n4 0.272055
R6869 VDD.n36 VDD.n35 0.272055
R6870 VDD.n47 VDD.n39 0.272055
R6871 VDD.n135 VDD.n134 0.2705
R6872 VDD.n22 VDD.n21 0.242579
R6873 VDD.n196 VDD.n185 0.239643
R6874 VDD.n368 VDD.n367 0.21542
R6875 VDD.n369 VDD.n368 0.18923
R6876 VDD.n415 VDD.n414 0.181952
R6877 VDD.n7 VDD.n5 0.17077
R6878 VDD.n33 VDD.n7 0.17077
R6879 VDD.n8 VDD.n6 0.17077
R6880 VDD.n33 VDD.n6 0.17077
R6881 VDD.n42 VDD.n41 0.17077
R6882 VDD.n45 VDD.n41 0.17077
R6883 VDD.n40 VDD.n2 0.17077
R6884 VDD.n45 VDD.n40 0.17077
R6885 VDD.n105 VDD.n104 0.149678
R6886 VDD.n205 VDD.n204 0.149643
R6887 VDD.n204 VDD.n202 0.149643
R6888 VDD.n415 VDD.n413 0.146702
R6889 VDD.n132 VDD.n131 0.142281
R6890 VDD.n104 VDD.n103 0.131185
R6891 VDD.n206 VDD.n201 0.127143
R6892 VDD.n158 VDD.n157 0.126253
R6893 VDD.n136 VDD.n135 0.120089
R6894 VDD.n195 VDD.n194 0.120071
R6895 VDD.n29 VDD.n28 0.11975
R6896 VDD.n28 VDD.n27 0.11975
R6897 VDD.n27 VDD.n11 0.11975
R6898 VDD.n23 VDD.n11 0.11975
R6899 VDD.n30 VDD.n10 0.11975
R6900 VDD.n26 VDD.n10 0.11975
R6901 VDD.n26 VDD.n25 0.11975
R6902 VDD.n25 VDD.n24 0.11975
R6903 VDD.n54 VDD.n53 0.11975
R6904 VDD.n53 VDD.n52 0.11975
R6905 VDD.n52 VDD.n3 0.11975
R6906 VDD.n48 VDD.n3 0.11975
R6907 VDD.n55 VDD.n1 0.11975
R6908 VDD.n51 VDD.n1 0.11975
R6909 VDD.n51 VDD.n50 0.11975
R6910 VDD.n50 VDD.n49 0.11975
R6911 VDD.n156 VDD.n155 0.115158
R6912 VDD.n137 VDD.n136 0.113925
R6913 VDD.n107 VDD.n106 0.113925
R6914 VDD.n133 VDD.n132 0.10776
R6915 VDD.n100 VDD.n99 0.106527
R6916 VDD.n240 VDD.n236 0.105016
R6917 VDD.n251 VDD.n236 0.105016
R6918 VDD.n253 VDD.n251 0.105016
R6919 VDD.n253 VDD.n252 0.105016
R6920 VDD.n252 VDD.n228 0.105016
R6921 VDD.n265 VDD.n228 0.105016
R6922 VDD.n267 VDD.n265 0.105016
R6923 VDD.n267 VDD.n266 0.105016
R6924 VDD.n266 VDD.n220 0.105016
R6925 VDD.n279 VDD.n220 0.105016
R6926 VDD.n282 VDD.n279 0.105016
R6927 VDD.n282 VDD.n281 0.105016
R6928 VDD.n281 VDD.n210 0.105016
R6929 VDD.n294 VDD.n210 0.105016
R6930 VDD.n172 VDD.n171 0.103753
R6931 VDD.n78 VDD.n77 0.101558
R6932 VDD.n102 VDD.n101 0.100363
R6933 VDD.n71 VDD.n70 0.0935717
R6934 VDD.n109 VDD.n108 0.0929658
R6935 VDD.n366 VDD.n365 0.0921268
R6936 VDD.n165 VDD.n164 0.0920411
R6937 VDD.n65 VDD.n64 0.0874283
R6938 VDD.n161 VDD.n160 0.080637
R6939 VDD.n67 VDD.n66 0.0791348
R6940 VDD.n112 VDD.n111 0.0757055
R6941 VDD.n63 VDD.n62 0.0751416
R6942 VDD.n111 VDD.n110 0.0744726
R6943 VDD.n174 VDD.n173 0.0723151
R6944 VDD.n169 VDD.n168 0.0692329
R6945 VDD.n368 VDD.n209 0.0672195
R6946 VDD.n75 VDD.n74 0.0671553
R6947 VDD.n108 VDD.n107 0.0646096
R6948 VDD.n62 VDD.n61 0.0634693
R6949 VDD.n138 VDD.n137 0.0624521
R6950 VDD.n114 VDD.n113 0.0624521
R6951 VDD.n69 VDD.n58 0.0622406
R6952 VDD.n31 VDD.n30 0.060125
R6953 VDD.n48 VDD.n47 0.060125
R6954 VDD.n49 VDD.n38 0.060125
R6955 VDD.n66 VDD.n65 0.0594761
R6956 VDD.n68 VDD.n67 0.0594761
R6957 VDD.n74 VDD.n73 0.0591689
R6958 VDD.n153 VDD.n152 0.0584452
R6959 VDD.n160 VDD.n159 0.0584452
R6960 VDD.n162 VDD.n161 0.0584452
R6961 VDD.n80 VDD.n68 0.0582474
R6962 VDD.n168 VDD.n167 0.0575205
R6963 VDD.n130 VDD.n129 0.0559795
R6964 VDD.n364 VDD.n310 0.0546935
R6965 VDD.n363 VDD.n295 0.0546935
R6966 VDD.n312 VDD.n309 0.0546935
R6967 VDD.n357 VDD.n296 0.0546935
R6968 VDD.n355 VDD.n308 0.0546935
R6969 VDD.n317 VDD.n297 0.0546935
R6970 VDD.n315 VDD.n307 0.0546935
R6971 VDD.n347 VDD.n298 0.0546935
R6972 VDD.n345 VDD.n306 0.0546935
R6973 VDD.n321 VDD.n299 0.0546935
R6974 VDD.n319 VDD.n305 0.0546935
R6975 VDD.n337 VDD.n300 0.0546935
R6976 VDD.n335 VDD.n304 0.0546935
R6977 VDD.n325 VDD.n301 0.0546935
R6978 VDD.n323 VDD.n303 0.0546935
R6979 VDD.n327 VDD.n302 0.0546935
R6980 VDD.n242 VDD.n241 0.0527581
R6981 VDD.n241 VDD.n239 0.0527581
R6982 VDD.n239 VDD.n237 0.0527581
R6983 VDD.n247 VDD.n237 0.0527581
R6984 VDD.n248 VDD.n247 0.0527581
R6985 VDD.n249 VDD.n248 0.0527581
R6986 VDD.n250 VDD.n249 0.0527581
R6987 VDD.n255 VDD.n254 0.0527581
R6988 VDD.n254 VDD.n235 0.0527581
R6989 VDD.n235 VDD.n229 0.0527581
R6990 VDD.n261 VDD.n229 0.0527581
R6991 VDD.n262 VDD.n261 0.0527581
R6992 VDD.n263 VDD.n262 0.0527581
R6993 VDD.n264 VDD.n263 0.0527581
R6994 VDD.n269 VDD.n268 0.0527581
R6995 VDD.n268 VDD.n227 0.0527581
R6996 VDD.n227 VDD.n221 0.0527581
R6997 VDD.n275 VDD.n221 0.0527581
R6998 VDD.n276 VDD.n275 0.0527581
R6999 VDD.n277 VDD.n276 0.0527581
R7000 VDD.n278 VDD.n277 0.0527581
R7001 VDD.n284 VDD.n283 0.0527581
R7002 VDD.n283 VDD.n219 0.0527581
R7003 VDD.n280 VDD.n219 0.0527581
R7004 VDD.n280 VDD.n214 0.0527581
R7005 VDD.n214 VDD.n213 0.0527581
R7006 VDD.n213 VDD.n211 0.0527581
R7007 VDD.n293 VDD.n211 0.0527581
R7008 VDD.n293 VDD.n292 0.0527581
R7009 VDD.n197 VDD.n195 0.0519286
R7010 VDD.n197 VDD.n196 0.0519286
R7011 VDD.n200 VDD.n185 0.0519286
R7012 VDD.n201 VDD.n200 0.0519286
R7013 VDD.n206 VDD.n205 0.0519286
R7014 VDD.n64 VDD.n63 0.0511826
R7015 VDD.n364 VDD.n363 0.0508226
R7016 VDD.n312 VDD.n295 0.0508226
R7017 VDD.n357 VDD.n309 0.0508226
R7018 VDD.n317 VDD.n308 0.0508226
R7019 VDD.n315 VDD.n297 0.0508226
R7020 VDD.n347 VDD.n307 0.0508226
R7021 VDD.n321 VDD.n306 0.0508226
R7022 VDD.n319 VDD.n299 0.0508226
R7023 VDD.n337 VDD.n305 0.0508226
R7024 VDD.n325 VDD.n304 0.0508226
R7025 VDD.n323 VDD.n301 0.0508226
R7026 VDD.n327 VDD.n303 0.0508226
R7027 VDD.n326 VDD.n302 0.0508226
R7028 VDD.n154 VDD.n153 0.0501233
R7029 VDD.n167 VDD.n166 0.0473493
R7030 VDD.n170 VDD.n169 0.0473493
R7031 VDD.n76 VDD.n75 0.0471894
R7032 VDD.n73 VDD.n72 0.0471894
R7033 VDD.n164 VDD.n163 0.0470411
R7034 VDD.n110 VDD.n109 0.0461164
R7035 VDD.n141 VDD.n140 0.0456716
R7036 VDD.n117 VDD.n116 0.0456716
R7037 VDD.n70 VDD.n69 0.0450393
R7038 VDD.n61 VDD.n60 0.0447321
R7039 VDD.n189 VDD.n183 0.0441954
R7040 VDD.n250 VDD.n234 0.0421129
R7041 VDD.n264 VDD.n226 0.0421129
R7042 VDD.n278 VDD.n218 0.0421129
R7043 VDD.n354 VDD.n296 0.0401774
R7044 VDD.n344 VDD.n298 0.0401774
R7045 VDD.n334 VDD.n300 0.0401774
R7046 VDD.n101 VDD.n100 0.0387192
R7047 VDD.n113 VDD.n112 0.0387192
R7048 VDD.n79 VDD.n78 0.0370529
R7049 VDD.n173 VDD.n172 0.0353288
R7050 VDD.n166 VDD.n165 0.0347123
R7051 VDD.n178 VDD.n176 0.0331712
R7052 VDD.n72 VDD.n71 0.0327526
R7053 VDD.n99 VDD.n98 0.0325548
R7054 VDD.n175 VDD.n174 0.0322466
R7055 VDD.n139 VDD.n138 0.0322466
R7056 VDD.n115 VDD.n114 0.0322466
R7057 VDD.n82 VDD.n58 0.0321382
R7058 VDD.n83 VDD.n82 0.0318362
R7059 VDD.n188 VDD.n187 0.0265682
R7060 VDD.n187 VDD.n186 0.0265682
R7061 VDD.n106 VDD.n105 0.0251575
R7062 VDD.n77 VDD.n76 0.0247662
R7063 VDD.n410 VDD.n409 0.024117
R7064 VDD.n403 VDD.n402 0.024117
R7065 VDD.n396 VDD.n395 0.024117
R7066 VDD.n389 VDD.n388 0.024117
R7067 VDD.n382 VDD.n381 0.024117
R7068 VDD.n375 VDD.n374 0.024117
R7069 VDD.n177 VDD.n145 0.0239247
R7070 VDD.n98 VDD.n97 0.0239247
R7071 VDD.n410 VDD.n405 0.0237979
R7072 VDD.n403 VDD.n398 0.0237979
R7073 VDD.n396 VDD.n391 0.0237979
R7074 VDD.n389 VDD.n384 0.0237979
R7075 VDD.n382 VDD.n377 0.0237979
R7076 VDD.n375 VDD.n370 0.0237979
R7077 VDD.n171 VDD.n170 0.023
R7078 VDD.n80 VDD.n79 0.0213874
R7079 VDD.n407 VDD.n406 0.020375
R7080 VDD.n408 VDD.n407 0.020375
R7081 VDD.n400 VDD.n399 0.020375
R7082 VDD.n401 VDD.n400 0.020375
R7083 VDD.n393 VDD.n392 0.020375
R7084 VDD.n394 VDD.n393 0.020375
R7085 VDD.n386 VDD.n385 0.020375
R7086 VDD.n387 VDD.n386 0.020375
R7087 VDD.n379 VDD.n378 0.020375
R7088 VDD.n380 VDD.n379 0.020375
R7089 VDD.n372 VDD.n371 0.020375
R7090 VDD.n373 VDD.n372 0.020375
R7091 VDD.n180 VDD.n144 0.0168356
R7092 VDD.n180 VDD.n179 0.0168356
R7093 VDD.n142 VDD.n119 0.0168356
R7094 VDD.n118 VDD.n84 0.0168356
R7095 VDD.n155 VDD.n154 0.0115959
R7096 VDD.n157 VDD.n156 0.0115959
R7097 VDD.n163 VDD.n162 0.0115959
R7098 VDD.n255 VDD.n234 0.0111452
R7099 VDD.n269 VDD.n226 0.0111452
R7100 VDD.n284 VDD.n218 0.0111452
R7101 VDD.n355 VDD.n354 0.0111452
R7102 VDD.n345 VDD.n344 0.0111452
R7103 VDD.n335 VDD.n334 0.0111452
R7104 VDD.n159 VDD.n158 0.0100548
R7105 VDD.n103 VDD.n102 0.00789726
R7106 VDD.n209 VDD.n184 0.00522745
R7107 VDD.n184 VDD.n57 0.00522745
R7108 VDD.n131 VDD.n130 0.00296575
R7109 VDD.n190 VDD.n189 0.00244773
R7110 VDD.n190 VDD.n0 0.00244773
R7111 VDD.n176 VDD.n175 0.00142466
R7112 VDD.n178 VDD.n177 0.00142466
R7113 VDD.n140 VDD.n139 0.00142466
R7114 VDD.n116 VDD.n115 0.00142466
R7115 F6.n6 F6.n5 7.13263
R7116 F6.n6 F6.n4 6.43746
R7117 F6.n12 F6.n1 6.43746
R7118 F6.n11 F6.n3 6.43746
R7119 F6.n5 F6.t9 3.8098
R7120 F6.n5 F6.t10 3.8098
R7121 F6.n4 F6.t13 3.8098
R7122 F6.n4 F6.t15 3.8098
R7123 F6.n1 F6.t11 3.8098
R7124 F6.n1 F6.t12 3.8098
R7125 F6.n3 F6.t14 3.8098
R7126 F6.n3 F6.t8 3.8098
R7127 F6.n9 F6.n8 3.34593
R7128 F6.n9 F6.n7 2.71593
R7129 F6.n12 F6.n0 2.71593
R7130 F6.n11 F6.n2 2.71593
R7131 F6.n7 F6.t0 2.06607
R7132 F6.n7 F6.t5 2.06607
R7133 F6.n8 F6.t3 2.06607
R7134 F6.n8 F6.t1 2.06607
R7135 F6.n0 F6.t6 2.06607
R7136 F6.n0 F6.t4 2.06607
R7137 F6.n2 F6.t2 2.06607
R7138 F6.n2 F6.t7 2.06607
R7139 F6.n10 F6.n6 0.382224
R7140 F6.n10 F6.n9 0.346437
R7141 F6.n12 F6.n11 0.138582
R7142 F6.n11 F6.n10 0.0627603
R7143 F6 F6.n12 0.00173288
R7144 OUT.n168 OUT.t3 29.4935
R7145 OUT.n61 OUT.n60 11.0705
R7146 OUT.n61 OUT.n59 11.0705
R7147 OUT.n67 OUT.n57 4.5005
R7148 OUT.n63 OUT.n57 4.5005
R7149 OUT.n67 OUT.n53 4.5005
R7150 OUT.n67 OUT.n66 4.5005
R7151 OUT.n66 OUT.n65 4.5005
R7152 OUT.n56 OUT.n54 4.27695
R7153 OUT.n56 OUT.n55 4.27695
R7154 OUT.n65 OUT.n62 2.24438
R7155 OUT.n63 OUT.n58 2.24438
R7156 OUT.n60 OUT.t2 1.6385
R7157 OUT.n60 OUT.t8 1.6385
R7158 OUT.n59 OUT.t1 1.6385
R7159 OUT.n59 OUT.t0 1.6385
R7160 OUT.n64 OUT.n50 1.51491
R7161 OUT.n70 OUT.n69 1.5005
R7162 OUT.n71 OUT.n49 1.5005
R7163 OUT.n73 OUT.n72 1.5005
R7164 OUT.n47 OUT.n46 1.5005
R7165 OUT.n78 OUT.n77 1.5005
R7166 OUT.n79 OUT.n45 1.5005
R7167 OUT.n81 OUT.n80 1.5005
R7168 OUT.n43 OUT.n42 1.5005
R7169 OUT.n86 OUT.n85 1.5005
R7170 OUT.n87 OUT.n41 1.5005
R7171 OUT.n89 OUT.n88 1.5005
R7172 OUT.n39 OUT.n38 1.5005
R7173 OUT.n94 OUT.n93 1.5005
R7174 OUT.n95 OUT.n37 1.5005
R7175 OUT.n97 OUT.n96 1.5005
R7176 OUT.n35 OUT.n34 1.5005
R7177 OUT.n102 OUT.n101 1.5005
R7178 OUT.n103 OUT.n33 1.5005
R7179 OUT.n105 OUT.n104 1.5005
R7180 OUT.n31 OUT.n30 1.5005
R7181 OUT.n110 OUT.n109 1.5005
R7182 OUT.n111 OUT.n29 1.5005
R7183 OUT.n113 OUT.n112 1.5005
R7184 OUT.n27 OUT.n26 1.5005
R7185 OUT.n118 OUT.n117 1.5005
R7186 OUT.n119 OUT.n25 1.5005
R7187 OUT.n121 OUT.n120 1.5005
R7188 OUT.n23 OUT.n22 1.5005
R7189 OUT.n126 OUT.n125 1.5005
R7190 OUT.n127 OUT.n21 1.5005
R7191 OUT.n129 OUT.n128 1.5005
R7192 OUT.n19 OUT.n18 1.5005
R7193 OUT.n134 OUT.n133 1.5005
R7194 OUT.n135 OUT.n17 1.5005
R7195 OUT.n137 OUT.n136 1.5005
R7196 OUT.n15 OUT.n14 1.5005
R7197 OUT.n142 OUT.n141 1.5005
R7198 OUT.n143 OUT.n13 1.5005
R7199 OUT.n145 OUT.n144 1.5005
R7200 OUT.n11 OUT.n10 1.5005
R7201 OUT.n150 OUT.n149 1.5005
R7202 OUT.n151 OUT.n9 1.5005
R7203 OUT.n153 OUT.n152 1.5005
R7204 OUT.n7 OUT.n6 1.5005
R7205 OUT.n158 OUT.n157 1.5005
R7206 OUT.n159 OUT.n5 1.5005
R7207 OUT.n161 OUT.n160 1.5005
R7208 OUT.n3 OUT.n2 1.5005
R7209 OUT.n166 OUT.n165 1.5005
R7210 OUT.n167 OUT.n1 1.5005
R7211 OUT.n173 OUT.n172 1.5005
R7212 OUT.n52 OUT.n51 1.5005
R7213 OUT.n69 OUT.n68 1.5005
R7214 OUT.n49 OUT.n48 1.5005
R7215 OUT.n74 OUT.n73 1.5005
R7216 OUT.n75 OUT.n47 1.5005
R7217 OUT.n77 OUT.n76 1.5005
R7218 OUT.n45 OUT.n44 1.5005
R7219 OUT.n82 OUT.n81 1.5005
R7220 OUT.n83 OUT.n43 1.5005
R7221 OUT.n85 OUT.n84 1.5005
R7222 OUT.n41 OUT.n40 1.5005
R7223 OUT.n90 OUT.n89 1.5005
R7224 OUT.n91 OUT.n39 1.5005
R7225 OUT.n93 OUT.n92 1.5005
R7226 OUT.n37 OUT.n36 1.5005
R7227 OUT.n98 OUT.n97 1.5005
R7228 OUT.n99 OUT.n35 1.5005
R7229 OUT.n101 OUT.n100 1.5005
R7230 OUT.n33 OUT.n32 1.5005
R7231 OUT.n106 OUT.n105 1.5005
R7232 OUT.n107 OUT.n31 1.5005
R7233 OUT.n109 OUT.n108 1.5005
R7234 OUT.n29 OUT.n28 1.5005
R7235 OUT.n114 OUT.n113 1.5005
R7236 OUT.n115 OUT.n27 1.5005
R7237 OUT.n117 OUT.n116 1.5005
R7238 OUT.n25 OUT.n24 1.5005
R7239 OUT.n122 OUT.n121 1.5005
R7240 OUT.n123 OUT.n23 1.5005
R7241 OUT.n125 OUT.n124 1.5005
R7242 OUT.n21 OUT.n20 1.5005
R7243 OUT.n130 OUT.n129 1.5005
R7244 OUT.n131 OUT.n19 1.5005
R7245 OUT.n133 OUT.n132 1.5005
R7246 OUT.n17 OUT.n16 1.5005
R7247 OUT.n138 OUT.n137 1.5005
R7248 OUT.n139 OUT.n15 1.5005
R7249 OUT.n141 OUT.n140 1.5005
R7250 OUT.n13 OUT.n12 1.5005
R7251 OUT.n146 OUT.n145 1.5005
R7252 OUT.n147 OUT.n11 1.5005
R7253 OUT.n149 OUT.n148 1.5005
R7254 OUT.n9 OUT.n8 1.5005
R7255 OUT.n154 OUT.n153 1.5005
R7256 OUT.n155 OUT.n7 1.5005
R7257 OUT.n157 OUT.n156 1.5005
R7258 OUT.n5 OUT.n4 1.5005
R7259 OUT.n162 OUT.n161 1.5005
R7260 OUT.n163 OUT.n3 1.5005
R7261 OUT.n165 OUT.n164 1.5005
R7262 OUT.n1 OUT.n0 1.5005
R7263 OUT.n174 OUT.n173 1.5005
R7264 OUT.n55 OUT.t4 0.9105
R7265 OUT.n55 OUT.t5 0.9105
R7266 OUT.n54 OUT.t7 0.9105
R7267 OUT.n54 OUT.t6 0.9105
R7268 OUT.n70 OUT.n50 0.76731
R7269 OUT.n172 OUT.n171 0.0668615
R7270 OUT.n69 OUT.n51 0.0284
R7271 OUT.n69 OUT.n49 0.0284
R7272 OUT.n73 OUT.n49 0.0284
R7273 OUT.n73 OUT.n47 0.0284
R7274 OUT.n77 OUT.n47 0.0284
R7275 OUT.n77 OUT.n45 0.0284
R7276 OUT.n81 OUT.n45 0.0284
R7277 OUT.n81 OUT.n43 0.0284
R7278 OUT.n85 OUT.n43 0.0284
R7279 OUT.n85 OUT.n41 0.0284
R7280 OUT.n89 OUT.n41 0.0284
R7281 OUT.n89 OUT.n39 0.0284
R7282 OUT.n93 OUT.n39 0.0284
R7283 OUT.n93 OUT.n37 0.0284
R7284 OUT.n97 OUT.n37 0.0284
R7285 OUT.n97 OUT.n35 0.0284
R7286 OUT.n101 OUT.n35 0.0284
R7287 OUT.n101 OUT.n33 0.0284
R7288 OUT.n105 OUT.n33 0.0284
R7289 OUT.n105 OUT.n31 0.0284
R7290 OUT.n109 OUT.n31 0.0284
R7291 OUT.n109 OUT.n29 0.0284
R7292 OUT.n113 OUT.n29 0.0284
R7293 OUT.n113 OUT.n27 0.0284
R7294 OUT.n117 OUT.n27 0.0284
R7295 OUT.n117 OUT.n25 0.0284
R7296 OUT.n121 OUT.n25 0.0284
R7297 OUT.n121 OUT.n23 0.0284
R7298 OUT.n125 OUT.n23 0.0284
R7299 OUT.n125 OUT.n21 0.0284
R7300 OUT.n129 OUT.n21 0.0284
R7301 OUT.n129 OUT.n19 0.0284
R7302 OUT.n133 OUT.n19 0.0284
R7303 OUT.n133 OUT.n17 0.0284
R7304 OUT.n137 OUT.n17 0.0284
R7305 OUT.n137 OUT.n15 0.0284
R7306 OUT.n141 OUT.n15 0.0284
R7307 OUT.n141 OUT.n13 0.0284
R7308 OUT.n145 OUT.n13 0.0284
R7309 OUT.n145 OUT.n11 0.0284
R7310 OUT.n149 OUT.n11 0.0284
R7311 OUT.n149 OUT.n9 0.0284
R7312 OUT.n153 OUT.n9 0.0284
R7313 OUT.n153 OUT.n7 0.0284
R7314 OUT.n157 OUT.n7 0.0284
R7315 OUT.n157 OUT.n5 0.0284
R7316 OUT.n161 OUT.n5 0.0284
R7317 OUT.n161 OUT.n3 0.0284
R7318 OUT.n165 OUT.n3 0.0284
R7319 OUT.n165 OUT.n1 0.0284
R7320 OUT.n173 OUT.n1 0.0284
R7321 OUT.n68 OUT.n48 0.0284
R7322 OUT.n74 OUT.n48 0.0284
R7323 OUT.n75 OUT.n74 0.0284
R7324 OUT.n76 OUT.n75 0.0284
R7325 OUT.n76 OUT.n44 0.0284
R7326 OUT.n82 OUT.n44 0.0284
R7327 OUT.n83 OUT.n82 0.0284
R7328 OUT.n84 OUT.n83 0.0284
R7329 OUT.n84 OUT.n40 0.0284
R7330 OUT.n90 OUT.n40 0.0284
R7331 OUT.n91 OUT.n90 0.0284
R7332 OUT.n92 OUT.n91 0.0284
R7333 OUT.n92 OUT.n36 0.0284
R7334 OUT.n98 OUT.n36 0.0284
R7335 OUT.n99 OUT.n98 0.0284
R7336 OUT.n100 OUT.n99 0.0284
R7337 OUT.n100 OUT.n32 0.0284
R7338 OUT.n106 OUT.n32 0.0284
R7339 OUT.n107 OUT.n106 0.0284
R7340 OUT.n108 OUT.n107 0.0284
R7341 OUT.n108 OUT.n28 0.0284
R7342 OUT.n114 OUT.n28 0.0284
R7343 OUT.n115 OUT.n114 0.0284
R7344 OUT.n116 OUT.n115 0.0284
R7345 OUT.n116 OUT.n24 0.0284
R7346 OUT.n122 OUT.n24 0.0284
R7347 OUT.n123 OUT.n122 0.0284
R7348 OUT.n124 OUT.n123 0.0284
R7349 OUT.n124 OUT.n20 0.0284
R7350 OUT.n130 OUT.n20 0.0284
R7351 OUT.n131 OUT.n130 0.0284
R7352 OUT.n132 OUT.n131 0.0284
R7353 OUT.n132 OUT.n16 0.0284
R7354 OUT.n138 OUT.n16 0.0284
R7355 OUT.n139 OUT.n138 0.0284
R7356 OUT.n140 OUT.n139 0.0284
R7357 OUT.n140 OUT.n12 0.0284
R7358 OUT.n146 OUT.n12 0.0284
R7359 OUT.n147 OUT.n146 0.0284
R7360 OUT.n148 OUT.n147 0.0284
R7361 OUT.n148 OUT.n8 0.0284
R7362 OUT.n154 OUT.n8 0.0284
R7363 OUT.n155 OUT.n154 0.0284
R7364 OUT.n156 OUT.n155 0.0284
R7365 OUT.n156 OUT.n4 0.0284
R7366 OUT.n162 OUT.n4 0.0284
R7367 OUT.n163 OUT.n162 0.0284
R7368 OUT.n164 OUT.n163 0.0284
R7369 OUT.n164 OUT.n0 0.0284
R7370 OUT.n174 OUT.n0 0.0284
R7371 OUT.n171 OUT.t19 0.0234592
R7372 OUT.n170 OUT.t14 0.0234592
R7373 OUT.n169 OUT.t10 0.0234592
R7374 OUT.n168 OUT.t20 0.0234592
R7375 OUT.n171 OUT.t13 0.0234592
R7376 OUT.n170 OUT.t12 0.0234592
R7377 OUT.n169 OUT.t9 0.0234592
R7378 OUT.n168 OUT.t18 0.0234592
R7379 OUT.n171 OUT.t17 0.0234592
R7380 OUT.n170 OUT.t16 0.0234592
R7381 OUT.n169 OUT.t15 0.0234592
R7382 OUT.n168 OUT.t11 0.0234592
R7383 OUT.n64 OUT.n63 0.023225
R7384 OUT.n67 OUT.n52 0.023225
R7385 OUT.n171 OUT.n170 0.0221244
R7386 OUT.n170 OUT.n169 0.0221244
R7387 OUT.n169 OUT.n168 0.0221244
R7388 OUT.n71 OUT.n70 0.0191
R7389 OUT.n72 OUT.n71 0.0191
R7390 OUT.n72 OUT.n46 0.0191
R7391 OUT.n78 OUT.n46 0.0191
R7392 OUT.n79 OUT.n78 0.0191
R7393 OUT.n80 OUT.n79 0.0191
R7394 OUT.n80 OUT.n42 0.0191
R7395 OUT.n86 OUT.n42 0.0191
R7396 OUT.n87 OUT.n86 0.0191
R7397 OUT.n88 OUT.n87 0.0191
R7398 OUT.n88 OUT.n38 0.0191
R7399 OUT.n94 OUT.n38 0.0191
R7400 OUT.n95 OUT.n94 0.0191
R7401 OUT.n96 OUT.n95 0.0191
R7402 OUT.n96 OUT.n34 0.0191
R7403 OUT.n102 OUT.n34 0.0191
R7404 OUT.n103 OUT.n102 0.0191
R7405 OUT.n104 OUT.n103 0.0191
R7406 OUT.n104 OUT.n30 0.0191
R7407 OUT.n110 OUT.n30 0.0191
R7408 OUT.n111 OUT.n110 0.0191
R7409 OUT.n112 OUT.n111 0.0191
R7410 OUT.n112 OUT.n26 0.0191
R7411 OUT.n118 OUT.n26 0.0191
R7412 OUT.n119 OUT.n118 0.0191
R7413 OUT.n120 OUT.n119 0.0191
R7414 OUT.n120 OUT.n22 0.0191
R7415 OUT.n126 OUT.n22 0.0191
R7416 OUT.n127 OUT.n126 0.0191
R7417 OUT.n128 OUT.n127 0.0191
R7418 OUT.n128 OUT.n18 0.0191
R7419 OUT.n134 OUT.n18 0.0191
R7420 OUT.n135 OUT.n134 0.0191
R7421 OUT.n136 OUT.n135 0.0191
R7422 OUT.n136 OUT.n14 0.0191
R7423 OUT.n142 OUT.n14 0.0191
R7424 OUT.n143 OUT.n142 0.0191
R7425 OUT.n144 OUT.n143 0.0191
R7426 OUT.n144 OUT.n10 0.0191
R7427 OUT.n150 OUT.n10 0.0191
R7428 OUT.n151 OUT.n150 0.0191
R7429 OUT.n152 OUT.n151 0.0191
R7430 OUT.n152 OUT.n6 0.0191
R7431 OUT.n158 OUT.n6 0.0191
R7432 OUT.n159 OUT.n158 0.0191
R7433 OUT.n160 OUT.n159 0.0191
R7434 OUT.n160 OUT.n2 0.0191
R7435 OUT.n166 OUT.n2 0.0191
R7436 OUT.n167 OUT.n166 0.0191
R7437 OUT.n172 OUT.n167 0.0191
R7438 OUT.n57 OUT.n56 0.0167857
R7439 OUT.n66 OUT.n61 0.0167857
R7440 OUT.n51 OUT.n50 0.0147371
R7441 OUT.n62 OUT.n53 0.0142466
R7442 OUT.n66 OUT.n58 0.0142466
R7443 OUT.n62 OUT.n57 0.0142466
R7444 OUT.n58 OUT.n53 0.0142466
R7445 OUT OUT.n174 0.0095
R7446 OUT.n65 OUT.n64 0.005675
R7447 OUT.n63 OUT.n52 0.005675
R7448 OUT.n68 OUT.n67 0.005675
R7449 a_5840_7613.t1 a_5840_7613.t0 25.621
R7450 a_22388_2038.t1 a_22388_2038.n1 21.2275
R7451 a_22388_2038.n1 a_22388_2038.t2 18.9805
R7452 a_22388_2038.n0 a_22388_2038.t5 17.5205
R7453 a_22388_2038.n0 a_22388_2038.t3 11.5588
R7454 a_22388_2038.n1 a_22388_2038.t4 11.4372
R7455 a_22388_2038.t1 a_22388_2038.t0 8.60523
R7456 a_22388_2038.t1 a_22388_2038.n0 8.27396
R7457 FREERUN.n75 FREERUN.t35 63.1691
R7458 FREERUN.t1 FREERUN.n26 58.6217
R7459 FREERUN.n9 FREERUN.t13 58.6217
R7460 FREERUN.n27 FREERUN.t1 55.3312
R7461 FREERUN.t13 FREERUN.n8 55.3312
R7462 FREERUN.n8 FREERUN.t14 39.8187
R7463 FREERUN.n9 FREERUN.t14 39.8187
R7464 FREERUN.n7 FREERUN.t32 39.8187
R7465 FREERUN.n10 FREERUN.t32 39.8187
R7466 FREERUN.n6 FREERUN.t5 39.8187
R7467 FREERUN.n11 FREERUN.t5 39.8187
R7468 FREERUN.n5 FREERUN.t24 39.8187
R7469 FREERUN.n12 FREERUN.t24 39.8187
R7470 FREERUN.n4 FREERUN.t9 39.8187
R7471 FREERUN.n13 FREERUN.t9 39.8187
R7472 FREERUN.n3 FREERUN.t27 39.8187
R7473 FREERUN.n14 FREERUN.t27 39.8187
R7474 FREERUN.n2 FREERUN.t15 39.8187
R7475 FREERUN.n15 FREERUN.t15 39.8187
R7476 FREERUN.n1 FREERUN.t3 39.8187
R7477 FREERUN.n16 FREERUN.t3 39.8187
R7478 FREERUN.t18 FREERUN.n0 39.8187
R7479 FREERUN.n17 FREERUN.t18 39.8187
R7480 FREERUN.n35 FREERUN.t37 39.8187
R7481 FREERUN.n18 FREERUN.t37 39.8187
R7482 FREERUN.n34 FREERUN.t23 39.8187
R7483 FREERUN.n19 FREERUN.t23 39.8187
R7484 FREERUN.n33 FREERUN.t40 39.8187
R7485 FREERUN.n20 FREERUN.t40 39.8187
R7486 FREERUN.n32 FREERUN.t30 39.8187
R7487 FREERUN.n21 FREERUN.t30 39.8187
R7488 FREERUN.n31 FREERUN.t4 39.8187
R7489 FREERUN.n22 FREERUN.t4 39.8187
R7490 FREERUN.n30 FREERUN.t34 39.8187
R7491 FREERUN.n23 FREERUN.t34 39.8187
R7492 FREERUN.n29 FREERUN.t7 39.8187
R7493 FREERUN.n24 FREERUN.t7 39.8187
R7494 FREERUN.n28 FREERUN.t25 39.8187
R7495 FREERUN.n25 FREERUN.t25 39.8187
R7496 FREERUN.n27 FREERUN.t12 39.8187
R7497 FREERUN.n26 FREERUN.t12 39.8187
R7498 FREERUN.n37 FREERUN.t38 37.0976
R7499 FREERUN.n47 FREERUN.t22 36.5005
R7500 FREERUN.t16 FREERUN.n64 36.5005
R7501 FREERUN.t22 FREERUN.n46 33.21
R7502 FREERUN.n65 FREERUN.t16 33.21
R7503 FREERUN.n48 FREERUN.n47 18.8035
R7504 FREERUN.n49 FREERUN.n48 18.8035
R7505 FREERUN.n50 FREERUN.n49 18.8035
R7506 FREERUN.n51 FREERUN.n50 18.8035
R7507 FREERUN.n52 FREERUN.n51 18.8035
R7508 FREERUN.n53 FREERUN.n52 18.8035
R7509 FREERUN.n54 FREERUN.n53 18.8035
R7510 FREERUN.n55 FREERUN.n54 18.8035
R7511 FREERUN.n56 FREERUN.n55 18.8035
R7512 FREERUN.n57 FREERUN.n56 18.8035
R7513 FREERUN.n58 FREERUN.n57 18.8035
R7514 FREERUN.n59 FREERUN.n58 18.8035
R7515 FREERUN.n60 FREERUN.n59 18.8035
R7516 FREERUN.n61 FREERUN.n60 18.8035
R7517 FREERUN.n62 FREERUN.n61 18.8035
R7518 FREERUN.n63 FREERUN.n62 18.8035
R7519 FREERUN.n64 FREERUN.n63 18.8035
R7520 FREERUN.n10 FREERUN.n9 18.8035
R7521 FREERUN.n11 FREERUN.n10 18.8035
R7522 FREERUN.n12 FREERUN.n11 18.8035
R7523 FREERUN.n13 FREERUN.n12 18.8035
R7524 FREERUN.n14 FREERUN.n13 18.8035
R7525 FREERUN.n15 FREERUN.n14 18.8035
R7526 FREERUN.n16 FREERUN.n15 18.8035
R7527 FREERUN.n17 FREERUN.n16 18.8035
R7528 FREERUN.n18 FREERUN.n17 18.8035
R7529 FREERUN.n19 FREERUN.n18 18.8035
R7530 FREERUN.n20 FREERUN.n19 18.8035
R7531 FREERUN.n21 FREERUN.n20 18.8035
R7532 FREERUN.n22 FREERUN.n21 18.8035
R7533 FREERUN.n23 FREERUN.n22 18.8035
R7534 FREERUN.n24 FREERUN.n23 18.8035
R7535 FREERUN.n25 FREERUN.n24 18.8035
R7536 FREERUN.n26 FREERUN.n25 18.8035
R7537 FREERUN.n65 FREERUN.t0 17.6975
R7538 FREERUN.n64 FREERUN.t0 17.6975
R7539 FREERUN.n66 FREERUN.t36 17.6975
R7540 FREERUN.n63 FREERUN.t36 17.6975
R7541 FREERUN.n67 FREERUN.t10 17.6975
R7542 FREERUN.n62 FREERUN.t10 17.6975
R7543 FREERUN.n68 FREERUN.t29 17.6975
R7544 FREERUN.n61 FREERUN.t29 17.6975
R7545 FREERUN.n69 FREERUN.t20 17.6975
R7546 FREERUN.n60 FREERUN.t20 17.6975
R7547 FREERUN.n70 FREERUN.t39 17.6975
R7548 FREERUN.n59 FREERUN.t39 17.6975
R7549 FREERUN.n71 FREERUN.t21 17.6975
R7550 FREERUN.n58 FREERUN.t21 17.6975
R7551 FREERUN.n72 FREERUN.t41 17.6975
R7552 FREERUN.n57 FREERUN.t41 17.6975
R7553 FREERUN.n73 FREERUN.t33 17.6975
R7554 FREERUN.n56 FREERUN.t33 17.6975
R7555 FREERUN.t8 FREERUN.n38 17.6975
R7556 FREERUN.n55 FREERUN.t8 17.6975
R7557 FREERUN.n39 FREERUN.t28 17.6975
R7558 FREERUN.n54 FREERUN.t28 17.6975
R7559 FREERUN.n40 FREERUN.t17 17.6975
R7560 FREERUN.n53 FREERUN.t17 17.6975
R7561 FREERUN.n41 FREERUN.t2 17.6975
R7562 FREERUN.n52 FREERUN.t2 17.6975
R7563 FREERUN.n42 FREERUN.t19 17.6975
R7564 FREERUN.n51 FREERUN.t19 17.6975
R7565 FREERUN.n43 FREERUN.t11 17.6975
R7566 FREERUN.n50 FREERUN.t11 17.6975
R7567 FREERUN.n44 FREERUN.t31 17.6975
R7568 FREERUN.n49 FREERUN.t31 17.6975
R7569 FREERUN.n45 FREERUN.t6 17.6975
R7570 FREERUN.n48 FREERUN.t6 17.6975
R7571 FREERUN.n46 FREERUN.t26 17.6975
R7572 FREERUN.n47 FREERUN.t26 17.6975
R7573 FREERUN.n46 FREERUN.n45 15.513
R7574 FREERUN.n45 FREERUN.n44 15.513
R7575 FREERUN.n44 FREERUN.n43 15.513
R7576 FREERUN.n43 FREERUN.n42 15.513
R7577 FREERUN.n42 FREERUN.n41 15.513
R7578 FREERUN.n41 FREERUN.n40 15.513
R7579 FREERUN.n40 FREERUN.n39 15.513
R7580 FREERUN.n39 FREERUN.n38 15.513
R7581 FREERUN.n73 FREERUN.n72 15.513
R7582 FREERUN.n72 FREERUN.n71 15.513
R7583 FREERUN.n71 FREERUN.n70 15.513
R7584 FREERUN.n70 FREERUN.n69 15.513
R7585 FREERUN.n69 FREERUN.n68 15.513
R7586 FREERUN.n68 FREERUN.n67 15.513
R7587 FREERUN.n67 FREERUN.n66 15.513
R7588 FREERUN.n66 FREERUN.n65 15.513
R7589 FREERUN.n8 FREERUN.n7 15.513
R7590 FREERUN.n7 FREERUN.n6 15.513
R7591 FREERUN.n6 FREERUN.n5 15.513
R7592 FREERUN.n5 FREERUN.n4 15.513
R7593 FREERUN.n4 FREERUN.n3 15.513
R7594 FREERUN.n3 FREERUN.n2 15.513
R7595 FREERUN.n2 FREERUN.n1 15.513
R7596 FREERUN.n1 FREERUN.n0 15.513
R7597 FREERUN.n35 FREERUN.n34 15.513
R7598 FREERUN.n34 FREERUN.n33 15.513
R7599 FREERUN.n33 FREERUN.n32 15.513
R7600 FREERUN.n32 FREERUN.n31 15.513
R7601 FREERUN.n31 FREERUN.n30 15.513
R7602 FREERUN.n30 FREERUN.n29 15.513
R7603 FREERUN.n29 FREERUN.n28 15.513
R7604 FREERUN.n28 FREERUN.n27 15.513
R7605 FREERUN.n74 FREERUN.n38 7.75675
R7606 FREERUN.n74 FREERUN.n73 7.75675
R7607 FREERUN.n36 FREERUN.n0 7.75675
R7608 FREERUN.n36 FREERUN.n35 7.75675
R7609 FREERUN.n37 FREERUN.n36 6.82995
R7610 FREERUN.n75 FREERUN.n74 6.82208
R7611 FREERUN FREERUN.n76 1.72963
R7612 FREERUN.n76 FREERUN.n75 0.77
R7613 FREERUN.n76 FREERUN.n37 0.487625
R7614 EX.n20 EX.n19 17.042
R7615 EX.n21 EX.n17 17.042
R7616 EX.n22 EX.n15 17.042
R7617 EX.n23 EX.n13 17.042
R7618 EX.n24 EX.n11 17.042
R7619 EX.n25 EX.n9 17.042
R7620 EX.n26 EX.n7 17.042
R7621 EX.n27 EX.n5 17.042
R7622 EX.n28 EX.n3 17.042
R7623 EX.n29 EX.n1 17.042
R7624 EX.n20 EX.n18 3.42767
R7625 EX.n21 EX.n16 3.42767
R7626 EX.n22 EX.n14 3.42767
R7627 EX.n23 EX.n12 3.42767
R7628 EX.n24 EX.n10 3.42767
R7629 EX.n25 EX.n8 3.42767
R7630 EX.n26 EX.n6 3.42767
R7631 EX.n27 EX.n4 3.42767
R7632 EX.n28 EX.n2 3.42767
R7633 EX.n29 EX.n0 3.42767
R7634 EX EX.n29 1.7762
R7635 EX.n19 EX.t10 1.6385
R7636 EX.n19 EX.t9 1.6385
R7637 EX.n17 EX.t1 1.6385
R7638 EX.n17 EX.t4 1.6385
R7639 EX.n15 EX.t12 1.6385
R7640 EX.n15 EX.t19 1.6385
R7641 EX.n13 EX.t16 1.6385
R7642 EX.n13 EX.t2 1.6385
R7643 EX.n11 EX.t8 1.6385
R7644 EX.n11 EX.t0 1.6385
R7645 EX.n9 EX.t7 1.6385
R7646 EX.n9 EX.t14 1.6385
R7647 EX.n7 EX.t11 1.6385
R7648 EX.n7 EX.t15 1.6385
R7649 EX.n5 EX.t18 1.6385
R7650 EX.n5 EX.t5 1.6385
R7651 EX.n3 EX.t13 1.6385
R7652 EX.n3 EX.t6 1.6385
R7653 EX.n1 EX.t17 1.6385
R7654 EX.n1 EX.t3 1.6385
R7655 EX.n18 EX.t30 0.607167
R7656 EX.n18 EX.t20 0.607167
R7657 EX.n16 EX.t34 0.607167
R7658 EX.n16 EX.t25 0.607167
R7659 EX.n14 EX.t23 0.607167
R7660 EX.n14 EX.t22 0.607167
R7661 EX.n12 EX.t29 0.607167
R7662 EX.n12 EX.t35 0.607167
R7663 EX.n10 EX.t21 0.607167
R7664 EX.n10 EX.t38 0.607167
R7665 EX.n8 EX.t27 0.607167
R7666 EX.n8 EX.t26 0.607167
R7667 EX.n6 EX.t24 0.607167
R7668 EX.n6 EX.t31 0.607167
R7669 EX.n4 EX.t37 0.607167
R7670 EX.n4 EX.t36 0.607167
R7671 EX.n2 EX.t39 0.607167
R7672 EX.n2 EX.t33 0.607167
R7673 EX.n0 EX.t32 0.607167
R7674 EX.n0 EX.t28 0.607167
R7675 EX.n21 EX.n20 0.1535
R7676 EX.n22 EX.n21 0.1535
R7677 EX.n23 EX.n22 0.1535
R7678 EX.n24 EX.n23 0.1535
R7679 EX.n25 EX.n24 0.1535
R7680 EX.n26 EX.n25 0.1535
R7681 EX.n27 EX.n26 0.1535
R7682 EX.n28 EX.n27 0.1535
R7683 EX.n29 EX.n28 0.1535
R7684 VCTRL VCTRL.t80 29.4036
R7685 VCTRL.n28 VCTRL.t8 14.1508
R7686 VCTRL.n18 VCTRL.t13 14.1508
R7687 VCTRL.n57 VCTRL.t67 14.1508
R7688 VCTRL.n47 VCTRL.t47 14.1508
R7689 VCTRL.n27 VCTRL.n1 11.5047
R7690 VCTRL.n26 VCTRL.n3 11.5047
R7691 VCTRL.n25 VCTRL.n5 11.5047
R7692 VCTRL.n24 VCTRL.n7 11.5047
R7693 VCTRL.n23 VCTRL.n9 11.5047
R7694 VCTRL.n22 VCTRL.n11 11.5047
R7695 VCTRL.n21 VCTRL.n13 11.5047
R7696 VCTRL.n20 VCTRL.n15 11.5047
R7697 VCTRL.n19 VCTRL.n17 11.5047
R7698 VCTRL.n56 VCTRL.n30 11.5047
R7699 VCTRL.n55 VCTRL.n32 11.5047
R7700 VCTRL.n54 VCTRL.n34 11.5047
R7701 VCTRL.n53 VCTRL.n36 11.5047
R7702 VCTRL.n52 VCTRL.n38 11.5047
R7703 VCTRL.n51 VCTRL.n40 11.5047
R7704 VCTRL.n50 VCTRL.n42 11.5047
R7705 VCTRL.n49 VCTRL.n44 11.5047
R7706 VCTRL.n48 VCTRL.n46 11.5047
R7707 VCTRL.n28 VCTRL.t66 4.19837
R7708 VCTRL.n18 VCTRL.t59 4.19837
R7709 VCTRL.n57 VCTRL.t24 4.19837
R7710 VCTRL.n47 VCTRL.t33 4.19837
R7711 VCTRL.n27 VCTRL.n0 3.21837
R7712 VCTRL.n26 VCTRL.n2 3.21837
R7713 VCTRL.n25 VCTRL.n4 3.21837
R7714 VCTRL.n24 VCTRL.n6 3.21837
R7715 VCTRL.n23 VCTRL.n8 3.21837
R7716 VCTRL.n22 VCTRL.n10 3.21837
R7717 VCTRL.n21 VCTRL.n12 3.21837
R7718 VCTRL.n20 VCTRL.n14 3.21837
R7719 VCTRL.n19 VCTRL.n16 3.21837
R7720 VCTRL.n56 VCTRL.n29 3.21837
R7721 VCTRL.n55 VCTRL.n31 3.21837
R7722 VCTRL.n54 VCTRL.n33 3.21837
R7723 VCTRL.n53 VCTRL.n35 3.21837
R7724 VCTRL.n52 VCTRL.n37 3.21837
R7725 VCTRL.n51 VCTRL.n39 3.21837
R7726 VCTRL.n50 VCTRL.n41 3.21837
R7727 VCTRL.n49 VCTRL.n43 3.21837
R7728 VCTRL.n48 VCTRL.n45 3.21837
R7729 VCTRL.n58 VCTRL.n28 1.73975
R7730 VCTRL.n1 VCTRL.t7 1.6385
R7731 VCTRL.n1 VCTRL.t17 1.6385
R7732 VCTRL.n3 VCTRL.t4 1.6385
R7733 VCTRL.n3 VCTRL.t14 1.6385
R7734 VCTRL.n5 VCTRL.t11 1.6385
R7735 VCTRL.n5 VCTRL.t18 1.6385
R7736 VCTRL.n7 VCTRL.t12 1.6385
R7737 VCTRL.n7 VCTRL.t6 1.6385
R7738 VCTRL.n9 VCTRL.t16 1.6385
R7739 VCTRL.n9 VCTRL.t3 1.6385
R7740 VCTRL.n11 VCTRL.t0 1.6385
R7741 VCTRL.n11 VCTRL.t9 1.6385
R7742 VCTRL.n13 VCTRL.t1 1.6385
R7743 VCTRL.n13 VCTRL.t10 1.6385
R7744 VCTRL.n15 VCTRL.t5 1.6385
R7745 VCTRL.n15 VCTRL.t15 1.6385
R7746 VCTRL.n17 VCTRL.t2 1.6385
R7747 VCTRL.n17 VCTRL.t19 1.6385
R7748 VCTRL.n30 VCTRL.t62 1.6385
R7749 VCTRL.n30 VCTRL.t61 1.6385
R7750 VCTRL.n32 VCTRL.t50 1.6385
R7751 VCTRL.n32 VCTRL.t42 1.6385
R7752 VCTRL.n34 VCTRL.t52 1.6385
R7753 VCTRL.n34 VCTRL.t70 1.6385
R7754 VCTRL.n36 VCTRL.t64 1.6385
R7755 VCTRL.n36 VCTRL.t48 1.6385
R7756 VCTRL.n38 VCTRL.t40 1.6385
R7757 VCTRL.n38 VCTRL.t54 1.6385
R7758 VCTRL.n40 VCTRL.t78 1.6385
R7759 VCTRL.n40 VCTRL.t55 1.6385
R7760 VCTRL.n42 VCTRL.t60 1.6385
R7761 VCTRL.n42 VCTRL.t49 1.6385
R7762 VCTRL.n44 VCTRL.t53 1.6385
R7763 VCTRL.n44 VCTRL.t51 1.6385
R7764 VCTRL.n46 VCTRL.t68 1.6385
R7765 VCTRL.n46 VCTRL.t65 1.6385
R7766 VCTRL.n0 VCTRL.t41 0.607167
R7767 VCTRL.n0 VCTRL.t73 0.607167
R7768 VCTRL.n2 VCTRL.t56 0.607167
R7769 VCTRL.n2 VCTRL.t45 0.607167
R7770 VCTRL.n4 VCTRL.t44 0.607167
R7771 VCTRL.n4 VCTRL.t63 0.607167
R7772 VCTRL.n6 VCTRL.t74 0.607167
R7773 VCTRL.n6 VCTRL.t43 0.607167
R7774 VCTRL.n8 VCTRL.t77 0.607167
R7775 VCTRL.n8 VCTRL.t58 0.607167
R7776 VCTRL.n10 VCTRL.t57 0.607167
R7777 VCTRL.n10 VCTRL.t46 0.607167
R7778 VCTRL.n12 VCTRL.t69 0.607167
R7779 VCTRL.n12 VCTRL.t76 0.607167
R7780 VCTRL.n14 VCTRL.t75 0.607167
R7781 VCTRL.n14 VCTRL.t79 0.607167
R7782 VCTRL.n16 VCTRL.t72 0.607167
R7783 VCTRL.n16 VCTRL.t71 0.607167
R7784 VCTRL.n29 VCTRL.t23 0.607167
R7785 VCTRL.n29 VCTRL.t35 0.607167
R7786 VCTRL.n31 VCTRL.t22 0.607167
R7787 VCTRL.n31 VCTRL.t28 0.607167
R7788 VCTRL.n33 VCTRL.t20 0.607167
R7789 VCTRL.n33 VCTRL.t26 0.607167
R7790 VCTRL.n35 VCTRL.t39 0.607167
R7791 VCTRL.n35 VCTRL.t32 0.607167
R7792 VCTRL.n37 VCTRL.t38 0.607167
R7793 VCTRL.n37 VCTRL.t30 0.607167
R7794 VCTRL.n39 VCTRL.t37 0.607167
R7795 VCTRL.n39 VCTRL.t29 0.607167
R7796 VCTRL.n41 VCTRL.t36 0.607167
R7797 VCTRL.n41 VCTRL.t31 0.607167
R7798 VCTRL.n43 VCTRL.t34 0.607167
R7799 VCTRL.n43 VCTRL.t21 0.607167
R7800 VCTRL.n45 VCTRL.t27 0.607167
R7801 VCTRL.n45 VCTRL.t25 0.607167
R7802 VCTRL VCTRL.n58 0.266975
R7803 VCTRL.n58 VCTRL.n57 0.21245
R7804 VCTRL.n28 VCTRL.n27 0.1679
R7805 VCTRL.n19 VCTRL.n18 0.1679
R7806 VCTRL.n57 VCTRL.n56 0.1679
R7807 VCTRL.n48 VCTRL.n47 0.1679
R7808 VCTRL.n27 VCTRL.n26 0.1535
R7809 VCTRL.n26 VCTRL.n25 0.1535
R7810 VCTRL.n25 VCTRL.n24 0.1535
R7811 VCTRL.n24 VCTRL.n23 0.1535
R7812 VCTRL.n23 VCTRL.n22 0.1535
R7813 VCTRL.n22 VCTRL.n21 0.1535
R7814 VCTRL.n21 VCTRL.n20 0.1535
R7815 VCTRL.n20 VCTRL.n19 0.1535
R7816 VCTRL.n56 VCTRL.n55 0.1535
R7817 VCTRL.n55 VCTRL.n54 0.1535
R7818 VCTRL.n54 VCTRL.n53 0.1535
R7819 VCTRL.n53 VCTRL.n52 0.1535
R7820 VCTRL.n52 VCTRL.n51 0.1535
R7821 VCTRL.n51 VCTRL.n50 0.1535
R7822 VCTRL.n50 VCTRL.n49 0.1535
R7823 VCTRL.n49 VCTRL.n48 0.1535
R7824 LF.n39 LF.n37 17.042
R7825 LF.n51 LF.n36 17.042
R7826 LF.n58 LF.n35 17.042
R7827 LF.n34 LF.n32 17.042
R7828 LF.n75 LF.n31 17.042
R7829 LF.n30 LF.n28 17.042
R7830 LF.n27 LF.n25 17.042
R7831 LF.n97 LF.n24 17.042
R7832 LF.n23 LF.n21 17.042
R7833 LF LF.n110 16.502
R7834 LF.n3 LF.t0 14.8576
R7835 LF.n104 LF.n103 4.5005
R7836 LF.n99 LF.n5 4.5005
R7837 LF.n6 LF.n5 4.5005
R7838 LF.n103 LF.n19 4.5005
R7839 LF.n99 LF.n19 4.5005
R7840 LF.n94 LF.n19 4.5005
R7841 LF.n92 LF.n19 4.5005
R7842 LF.n89 LF.n19 4.5005
R7843 LF.n87 LF.n19 4.5005
R7844 LF.n84 LF.n19 4.5005
R7845 LF.n82 LF.n19 4.5005
R7846 LF.n79 LF.n19 4.5005
R7847 LF.n77 LF.n19 4.5005
R7848 LF.n72 LF.n19 4.5005
R7849 LF.n70 LF.n19 4.5005
R7850 LF.n67 LF.n19 4.5005
R7851 LF.n65 LF.n19 4.5005
R7852 LF.n62 LF.n19 4.5005
R7853 LF.n60 LF.n19 4.5005
R7854 LF.n55 LF.n19 4.5005
R7855 LF.n53 LF.n19 4.5005
R7856 LF.n48 LF.n19 4.5005
R7857 LF.n46 LF.n19 4.5005
R7858 LF.n43 LF.n19 4.5005
R7859 LF.n41 LF.n19 4.5005
R7860 LF.n109 LF.n108 3.38042
R7861 LF.n39 LF.n38 3.38042
R7862 LF.n51 LF.n50 3.38042
R7863 LF.n58 LF.n57 3.38042
R7864 LF.n34 LF.n33 3.38042
R7865 LF.n75 LF.n74 3.38042
R7866 LF.n30 LF.n29 3.38042
R7867 LF.n27 LF.n26 3.38042
R7868 LF.n97 LF.n96 3.38042
R7869 LF.n23 LF.n22 3.38042
R7870 LF.n106 LF.n105 2.25041
R7871 LF.n100 LF.n18 2.25041
R7872 LF.n104 LF.n17 2.24525
R7873 LF.n104 LF.n16 2.24525
R7874 LF.n104 LF.n15 2.24525
R7875 LF.n104 LF.n14 2.24525
R7876 LF.n104 LF.n13 2.24525
R7877 LF.n104 LF.n12 2.24525
R7878 LF.n104 LF.n11 2.24525
R7879 LF.n104 LF.n10 2.24525
R7880 LF.n104 LF.n9 2.24525
R7881 LF.n104 LF.n8 2.24525
R7882 LF.n104 LF.n7 2.24525
R7883 LF.n20 LF.n5 2.24525
R7884 LF.n93 LF.n5 2.24525
R7885 LF.n88 LF.n5 2.24525
R7886 LF.n83 LF.n5 2.24525
R7887 LF.n78 LF.n5 2.24525
R7888 LF.n71 LF.n5 2.24525
R7889 LF.n66 LF.n5 2.24525
R7890 LF.n61 LF.n5 2.24525
R7891 LF.n54 LF.n5 2.24525
R7892 LF.n47 LF.n5 2.24525
R7893 LF.n42 LF.n5 2.24525
R7894 LF.n19 LF.n1 2.24525
R7895 LF.n110 LF.t36 1.6385
R7896 LF.n110 LF.t23 1.6385
R7897 LF.n37 LF.t27 1.6385
R7898 LF.n37 LF.t38 1.6385
R7899 LF.n36 LF.t25 1.6385
R7900 LF.n36 LF.t29 1.6385
R7901 LF.n35 LF.t31 1.6385
R7902 LF.n35 LF.t32 1.6385
R7903 LF.n32 LF.t30 1.6385
R7904 LF.n32 LF.t40 1.6385
R7905 LF.n31 LF.t24 1.6385
R7906 LF.n31 LF.t21 1.6385
R7907 LF.n28 LF.t39 1.6385
R7908 LF.n28 LF.t35 1.6385
R7909 LF.n25 LF.t22 1.6385
R7910 LF.n25 LF.t28 1.6385
R7911 LF.n24 LF.t33 1.6385
R7912 LF.n24 LF.t26 1.6385
R7913 LF.n21 LF.t37 1.6385
R7914 LF.n21 LF.t34 1.6385
R7915 LF.n103 LF.n102 1.5005
R7916 LF.n101 LF.n100 1.5005
R7917 LF.n99 LF.n98 1.5005
R7918 LF.n95 LF.n94 1.5005
R7919 LF.n92 LF.n91 1.5005
R7920 LF.n90 LF.n89 1.5005
R7921 LF.n87 LF.n86 1.5005
R7922 LF.n85 LF.n84 1.5005
R7923 LF.n82 LF.n81 1.5005
R7924 LF.n80 LF.n79 1.5005
R7925 LF.n77 LF.n76 1.5005
R7926 LF.n73 LF.n72 1.5005
R7927 LF.n70 LF.n69 1.5005
R7928 LF.n68 LF.n67 1.5005
R7929 LF.n65 LF.n64 1.5005
R7930 LF.n63 LF.n62 1.5005
R7931 LF.n60 LF.n59 1.5005
R7932 LF.n56 LF.n55 1.5005
R7933 LF.n53 LF.n52 1.5005
R7934 LF.n49 LF.n48 1.5005
R7935 LF.n46 LF.n45 1.5005
R7936 LF.n44 LF.n43 1.5005
R7937 LF.n41 LF.n40 1.5005
R7938 LF.n6 LF.n0 1.5005
R7939 LF.n107 LF.n106 1.5005
R7940 LF.n108 LF.t14 0.607167
R7941 LF.n108 LF.t20 0.607167
R7942 LF.n38 LF.t16 0.607167
R7943 LF.n38 LF.t7 0.607167
R7944 LF.n50 LF.t18 0.607167
R7945 LF.n50 LF.t3 0.607167
R7946 LF.n57 LF.t1 0.607167
R7947 LF.n57 LF.t5 0.607167
R7948 LF.n33 LF.t2 0.607167
R7949 LF.n33 LF.t9 0.607167
R7950 LF.n74 LF.t19 0.607167
R7951 LF.n74 LF.t10 0.607167
R7952 LF.n29 LF.t6 0.607167
R7953 LF.n29 LF.t11 0.607167
R7954 LF.n26 LF.t8 0.607167
R7955 LF.n26 LF.t15 0.607167
R7956 LF.n96 LF.t4 0.607167
R7957 LF.n96 LF.t17 0.607167
R7958 LF.n22 LF.t13 0.607167
R7959 LF.n22 LF.t12 0.607167
R7960 LF LF.n109 0.5405
R7961 LF.n5 LF.n4 0.119279
R7962 LF.n2 LF.t47 0.063
R7963 LF.n4 LF.t50 0.063
R7964 LF.n2 LF.t49 0.063
R7965 LF.n4 LF.t44 0.063
R7966 LF.n2 LF.t41 0.063
R7967 LF.n4 LF.t45 0.063
R7968 LF.n2 LF.t48 0.063
R7969 LF.n4 LF.t43 0.063
R7970 LF.n2 LF.t42 0.063
R7971 LF.n4 LF.t46 0.063
R7972 LF.n100 LF.n99 0.0235579
R7973 LF.n102 LF.n101 0.0235579
R7974 LF.n101 LF.n98 0.0235579
R7975 LF.n95 LF.n91 0.0235579
R7976 LF.n91 LF.n90 0.0235579
R7977 LF.n86 LF.n85 0.0235579
R7978 LF.n81 LF.n80 0.0235579
R7979 LF.n80 LF.n76 0.0235579
R7980 LF.n73 LF.n69 0.0235579
R7981 LF.n69 LF.n68 0.0235579
R7982 LF.n64 LF.n63 0.0235579
R7983 LF.n63 LF.n59 0.0235579
R7984 LF.n56 LF.n52 0.0235579
R7985 LF.n49 LF.n45 0.0235579
R7986 LF.n45 LF.n44 0.0235579
R7987 LF.n40 LF.n0 0.0235579
R7988 LF.n107 LF.n0 0.0235579
R7989 LF.n85 LF.n30 0.0209545
R7990 LF.n58 LF.n56 0.0209545
R7991 LF.n86 LF.n27 0.0202107
R7992 LF.n52 LF.n51 0.0202107
R7993 LF.n76 LF.n75 0.0150041
R7994 LF.n64 LF.n34 0.0150041
R7995 LF.n97 LF.n95 0.0142603
R7996 LF.n44 LF.n39 0.0142603
R7997 LF.n100 LF.n20 0.0124995
R7998 LF.n94 LF.n17 0.0124995
R7999 LF.n94 LF.n93 0.0124995
R8000 LF.n89 LF.n16 0.0124995
R8001 LF.n89 LF.n88 0.0124995
R8002 LF.n84 LF.n15 0.0124995
R8003 LF.n84 LF.n83 0.0124995
R8004 LF.n79 LF.n14 0.0124995
R8005 LF.n79 LF.n78 0.0124995
R8006 LF.n72 LF.n13 0.0124995
R8007 LF.n72 LF.n71 0.0124995
R8008 LF.n67 LF.n12 0.0124995
R8009 LF.n67 LF.n66 0.0124995
R8010 LF.n62 LF.n11 0.0124995
R8011 LF.n62 LF.n61 0.0124995
R8012 LF.n55 LF.n10 0.0124995
R8013 LF.n55 LF.n54 0.0124995
R8014 LF.n48 LF.n9 0.0124995
R8015 LF.n48 LF.n47 0.0124995
R8016 LF.n43 LF.n8 0.0124995
R8017 LF.n43 LF.n42 0.0124995
R8018 LF.n7 LF.n6 0.0124995
R8019 LF.n6 LF.n1 0.0124995
R8020 LF.n99 LF.n17 0.0124995
R8021 LF.n92 LF.n16 0.0124995
R8022 LF.n87 LF.n15 0.0124995
R8023 LF.n82 LF.n14 0.0124995
R8024 LF.n77 LF.n13 0.0124995
R8025 LF.n70 LF.n12 0.0124995
R8026 LF.n65 LF.n11 0.0124995
R8027 LF.n60 LF.n10 0.0124995
R8028 LF.n53 LF.n9 0.0124995
R8029 LF.n46 LF.n8 0.0124995
R8030 LF.n41 LF.n7 0.0124995
R8031 LF.n103 LF.n20 0.0124995
R8032 LF.n93 LF.n92 0.0124995
R8033 LF.n88 LF.n87 0.0124995
R8034 LF.n83 LF.n82 0.0124995
R8035 LF.n78 LF.n77 0.0124995
R8036 LF.n71 LF.n70 0.0124995
R8037 LF.n66 LF.n65 0.0124995
R8038 LF.n61 LF.n60 0.0124995
R8039 LF.n54 LF.n53 0.0124995
R8040 LF.n47 LF.n46 0.0124995
R8041 LF.n42 LF.n41 0.0124995
R8042 LF.n106 LF.n1 0.0124995
R8043 LF.n3 LF.n2 0.0109762
R8044 LF.n4 LF.n3 0.0109762
R8045 LF.n98 LF.n97 0.00979752
R8046 LF.n40 LF.n39 0.00979752
R8047 LF.n75 LF.n73 0.00905372
R8048 LF.n68 LF.n34 0.00905372
R8049 LF.n102 LF.n23 0.00830992
R8050 LF.n109 LF.n107 0.00830992
R8051 LF.n90 LF.n27 0.00384711
R8052 LF.n51 LF.n49 0.00384711
R8053 LF.n81 LF.n30 0.00310331
R8054 LF.n59 LF.n58 0.00310331
R8055 LF.n105 LF.n104 0.0021844
R8056 LF.n19 LF.n18 0.0021844
R8057 LF.n104 LF.n18 0.0021844
R8058 LF.n105 LF.n5 0.0021844
R8059 a_n558_2704.n3 a_n558_2704.t8 39.434
R8060 a_n558_2704.n0 a_n558_2704.t6 39.3425
R8061 a_n558_2704.n0 a_n558_2704.t7 29.4555
R8062 a_n558_2704.n3 a_n558_2704.t5 29.3205
R8063 a_n558_2704.n1 a_n558_2704.t4 28.7301
R8064 a_n558_2704.n1 a_n558_2704.t3 18.7615
R8065 a_n558_2704.n2 a_n558_2704.t1 13.7342
R8066 a_n558_2704.n1 a_n558_2704.t2 13.5055
R8067 a_n558_2704.n0 a_n558_2704.n1 9.0247
R8068 a_n558_2704.n2 a_n558_2704.n3 7.96025
R8069 a_n558_2704.t0 a_n558_2704.n2 6.3271
R8070 a_n558_2704.n2 a_n558_2704.n0 1.39825
R8071 a_n17351_68.t21 a_n17351_68.n64 58.6217
R8072 a_n17351_68.n47 a_n17351_68.t34 58.6217
R8073 a_n17351_68.n65 a_n17351_68.t21 55.3312
R8074 a_n17351_68.t34 a_n17351_68.n46 55.3312
R8075 a_n17351_68.n46 a_n17351_68.t12 39.8187
R8076 a_n17351_68.n47 a_n17351_68.t12 39.8187
R8077 a_n17351_68.n45 a_n17351_68.t8 39.8187
R8078 a_n17351_68.n48 a_n17351_68.t8 39.8187
R8079 a_n17351_68.n44 a_n17351_68.t3 39.8187
R8080 a_n17351_68.n49 a_n17351_68.t3 39.8187
R8081 a_n17351_68.n43 a_n17351_68.t40 39.8187
R8082 a_n17351_68.n50 a_n17351_68.t40 39.8187
R8083 a_n17351_68.n42 a_n17351_68.t39 39.8187
R8084 a_n17351_68.n51 a_n17351_68.t39 39.8187
R8085 a_n17351_68.n41 a_n17351_68.t37 39.8187
R8086 a_n17351_68.n52 a_n17351_68.t37 39.8187
R8087 a_n17351_68.n40 a_n17351_68.t15 39.8187
R8088 a_n17351_68.n53 a_n17351_68.t15 39.8187
R8089 a_n17351_68.n39 a_n17351_68.t14 39.8187
R8090 a_n17351_68.n54 a_n17351_68.t14 39.8187
R8091 a_n17351_68.t9 a_n17351_68.n38 39.8187
R8092 a_n17351_68.n55 a_n17351_68.t9 39.8187
R8093 a_n17351_68.n73 a_n17351_68.t5 39.8187
R8094 a_n17351_68.n56 a_n17351_68.t5 39.8187
R8095 a_n17351_68.n72 a_n17351_68.t4 39.8187
R8096 a_n17351_68.n57 a_n17351_68.t4 39.8187
R8097 a_n17351_68.n71 a_n17351_68.t41 39.8187
R8098 a_n17351_68.n58 a_n17351_68.t41 39.8187
R8099 a_n17351_68.n70 a_n17351_68.t19 39.8187
R8100 a_n17351_68.n59 a_n17351_68.t19 39.8187
R8101 a_n17351_68.n69 a_n17351_68.t17 39.8187
R8102 a_n17351_68.n60 a_n17351_68.t17 39.8187
R8103 a_n17351_68.n68 a_n17351_68.t16 39.8187
R8104 a_n17351_68.n61 a_n17351_68.t16 39.8187
R8105 a_n17351_68.n67 a_n17351_68.t11 39.8187
R8106 a_n17351_68.n62 a_n17351_68.t11 39.8187
R8107 a_n17351_68.n66 a_n17351_68.t7 39.8187
R8108 a_n17351_68.n63 a_n17351_68.t7 39.8187
R8109 a_n17351_68.n65 a_n17351_68.t6 39.8187
R8110 a_n17351_68.n64 a_n17351_68.t6 39.8187
R8111 a_n17351_68.n10 a_n17351_68.t35 36.5005
R8112 a_n17351_68.t27 a_n17351_68.n27 36.5005
R8113 a_n17351_68.t35 a_n17351_68.n9 33.21
R8114 a_n17351_68.n28 a_n17351_68.t27 33.21
R8115 a_n17351_68.n11 a_n17351_68.n10 18.8035
R8116 a_n17351_68.n12 a_n17351_68.n11 18.8035
R8117 a_n17351_68.n13 a_n17351_68.n12 18.8035
R8118 a_n17351_68.n14 a_n17351_68.n13 18.8035
R8119 a_n17351_68.n15 a_n17351_68.n14 18.8035
R8120 a_n17351_68.n16 a_n17351_68.n15 18.8035
R8121 a_n17351_68.n17 a_n17351_68.n16 18.8035
R8122 a_n17351_68.n18 a_n17351_68.n17 18.8035
R8123 a_n17351_68.n19 a_n17351_68.n18 18.8035
R8124 a_n17351_68.n20 a_n17351_68.n19 18.8035
R8125 a_n17351_68.n21 a_n17351_68.n20 18.8035
R8126 a_n17351_68.n22 a_n17351_68.n21 18.8035
R8127 a_n17351_68.n23 a_n17351_68.n22 18.8035
R8128 a_n17351_68.n24 a_n17351_68.n23 18.8035
R8129 a_n17351_68.n25 a_n17351_68.n24 18.8035
R8130 a_n17351_68.n26 a_n17351_68.n25 18.8035
R8131 a_n17351_68.n27 a_n17351_68.n26 18.8035
R8132 a_n17351_68.n48 a_n17351_68.n47 18.8035
R8133 a_n17351_68.n49 a_n17351_68.n48 18.8035
R8134 a_n17351_68.n50 a_n17351_68.n49 18.8035
R8135 a_n17351_68.n51 a_n17351_68.n50 18.8035
R8136 a_n17351_68.n52 a_n17351_68.n51 18.8035
R8137 a_n17351_68.n53 a_n17351_68.n52 18.8035
R8138 a_n17351_68.n54 a_n17351_68.n53 18.8035
R8139 a_n17351_68.n55 a_n17351_68.n54 18.8035
R8140 a_n17351_68.n56 a_n17351_68.n55 18.8035
R8141 a_n17351_68.n57 a_n17351_68.n56 18.8035
R8142 a_n17351_68.n58 a_n17351_68.n57 18.8035
R8143 a_n17351_68.n59 a_n17351_68.n58 18.8035
R8144 a_n17351_68.n60 a_n17351_68.n59 18.8035
R8145 a_n17351_68.n61 a_n17351_68.n60 18.8035
R8146 a_n17351_68.n62 a_n17351_68.n61 18.8035
R8147 a_n17351_68.n63 a_n17351_68.n62 18.8035
R8148 a_n17351_68.n64 a_n17351_68.n63 18.8035
R8149 a_n17351_68.n28 a_n17351_68.t33 17.6975
R8150 a_n17351_68.n27 a_n17351_68.t33 17.6975
R8151 a_n17351_68.n29 a_n17351_68.t18 17.6975
R8152 a_n17351_68.n26 a_n17351_68.t18 17.6975
R8153 a_n17351_68.n30 a_n17351_68.t31 17.6975
R8154 a_n17351_68.n25 a_n17351_68.t31 17.6975
R8155 a_n17351_68.n31 a_n17351_68.t24 17.6975
R8156 a_n17351_68.n24 a_n17351_68.t24 17.6975
R8157 a_n17351_68.n32 a_n17351_68.t29 17.6975
R8158 a_n17351_68.n23 a_n17351_68.t29 17.6975
R8159 a_n17351_68.n33 a_n17351_68.t22 17.6975
R8160 a_n17351_68.n22 a_n17351_68.t22 17.6975
R8161 a_n17351_68.n34 a_n17351_68.t26 17.6975
R8162 a_n17351_68.n21 a_n17351_68.t26 17.6975
R8163 a_n17351_68.n35 a_n17351_68.t10 17.6975
R8164 a_n17351_68.n20 a_n17351_68.t10 17.6975
R8165 a_n17351_68.n36 a_n17351_68.t25 17.6975
R8166 a_n17351_68.n19 a_n17351_68.t25 17.6975
R8167 a_n17351_68.t2 a_n17351_68.n1 17.6975
R8168 a_n17351_68.n18 a_n17351_68.t2 17.6975
R8169 a_n17351_68.n2 a_n17351_68.t28 17.6975
R8170 a_n17351_68.n17 a_n17351_68.t28 17.6975
R8171 a_n17351_68.n3 a_n17351_68.t38 17.6975
R8172 a_n17351_68.n16 a_n17351_68.t38 17.6975
R8173 a_n17351_68.n4 a_n17351_68.t20 17.6975
R8174 a_n17351_68.n15 a_n17351_68.t20 17.6975
R8175 a_n17351_68.n5 a_n17351_68.t32 17.6975
R8176 a_n17351_68.n14 a_n17351_68.t32 17.6975
R8177 a_n17351_68.n6 a_n17351_68.t13 17.6975
R8178 a_n17351_68.n13 a_n17351_68.t13 17.6975
R8179 a_n17351_68.n7 a_n17351_68.t30 17.6975
R8180 a_n17351_68.n12 a_n17351_68.t30 17.6975
R8181 a_n17351_68.n8 a_n17351_68.t23 17.6975
R8182 a_n17351_68.n11 a_n17351_68.t23 17.6975
R8183 a_n17351_68.n9 a_n17351_68.t36 17.6975
R8184 a_n17351_68.n10 a_n17351_68.t36 17.6975
R8185 a_n17351_68.n9 a_n17351_68.n8 15.513
R8186 a_n17351_68.n8 a_n17351_68.n7 15.513
R8187 a_n17351_68.n7 a_n17351_68.n6 15.513
R8188 a_n17351_68.n6 a_n17351_68.n5 15.513
R8189 a_n17351_68.n5 a_n17351_68.n4 15.513
R8190 a_n17351_68.n4 a_n17351_68.n3 15.513
R8191 a_n17351_68.n3 a_n17351_68.n2 15.513
R8192 a_n17351_68.n2 a_n17351_68.n1 15.513
R8193 a_n17351_68.n36 a_n17351_68.n35 15.513
R8194 a_n17351_68.n35 a_n17351_68.n34 15.513
R8195 a_n17351_68.n34 a_n17351_68.n33 15.513
R8196 a_n17351_68.n33 a_n17351_68.n32 15.513
R8197 a_n17351_68.n32 a_n17351_68.n31 15.513
R8198 a_n17351_68.n31 a_n17351_68.n30 15.513
R8199 a_n17351_68.n30 a_n17351_68.n29 15.513
R8200 a_n17351_68.n29 a_n17351_68.n28 15.513
R8201 a_n17351_68.n46 a_n17351_68.n45 15.513
R8202 a_n17351_68.n45 a_n17351_68.n44 15.513
R8203 a_n17351_68.n44 a_n17351_68.n43 15.513
R8204 a_n17351_68.n43 a_n17351_68.n42 15.513
R8205 a_n17351_68.n42 a_n17351_68.n41 15.513
R8206 a_n17351_68.n41 a_n17351_68.n40 15.513
R8207 a_n17351_68.n40 a_n17351_68.n39 15.513
R8208 a_n17351_68.n39 a_n17351_68.n38 15.513
R8209 a_n17351_68.n73 a_n17351_68.n72 15.513
R8210 a_n17351_68.n72 a_n17351_68.n71 15.513
R8211 a_n17351_68.n71 a_n17351_68.n70 15.513
R8212 a_n17351_68.n70 a_n17351_68.n69 15.513
R8213 a_n17351_68.n69 a_n17351_68.n68 15.513
R8214 a_n17351_68.n68 a_n17351_68.n67 15.513
R8215 a_n17351_68.n67 a_n17351_68.n66 15.513
R8216 a_n17351_68.n66 a_n17351_68.n65 15.513
R8217 a_n17351_68.n75 a_n17351_68.t1 14.2059
R8218 a_n17351_68.n37 a_n17351_68.n1 7.75675
R8219 a_n17351_68.n37 a_n17351_68.n36 7.75675
R8220 a_n17351_68.n74 a_n17351_68.n38 7.75675
R8221 a_n17351_68.n74 a_n17351_68.n73 7.75675
R8222 a_n17351_68.t0 a_n17351_68.n75 4.23734
R8223 a_n17351_68.n0 a_n17351_68.n37 0.633736
R8224 a_n17351_68.n0 a_n17351_68.n74 0.59343
R8225 a_n17351_68.n0 a_n17351_68.n75 2.39173
R8226 a_22203_n358.n5 a_22203_n358.t15 31.6987
R8227 a_22203_n358.n6 a_22203_n358.t17 18.6885
R8228 a_22203_n358.n7 a_22203_n358.t14 18.6885
R8229 a_22203_n358.n5 a_22203_n358.t18 18.6885
R8230 a_22203_n358.n10 a_22203_n358.t16 13.907
R8231 a_22203_n358.n9 a_22203_n358.t12 13.8462
R8232 a_22203_n358.n11 a_22203_n358.t20 13.8462
R8233 a_22203_n358.n9 a_22203_n358.t9 12.1185
R8234 a_22203_n358.n11 a_22203_n358.t19 12.1185
R8235 a_22203_n358.n10 a_22203_n358.t8 12.0455
R8236 a_22203_n358.n6 a_22203_n358.t10 11.1938
R8237 a_22203_n358.n7 a_22203_n358.t13 11.1938
R8238 a_22203_n358.n5 a_22203_n358.t11 11.1938
R8239 a_22203_n358.n1 a_22203_n358.n9 10.6383
R8240 a_22203_n358.n7 a_22203_n358.n6 10.5449
R8241 a_22203_n358.n1 a_22203_n358.n11 10.2813
R8242 a_22203_n358.n1 a_22203_n358.n10 10.2813
R8243 a_22203_n358.n0 a_22203_n358.n4 7.33746
R8244 a_22203_n358.n8 a_22203_n358.n5 6.48939
R8245 a_22203_n358.n0 a_22203_n358.n3 6.46093
R8246 a_22203_n358.n12 a_22203_n358.n0 6.01368
R8247 a_22203_n358.n0 a_22203_n358.n2 5.4118
R8248 a_22203_n358.n8 a_22203_n358.n7 4.05606
R8249 a_22203_n358.n4 a_22203_n358.t4 3.6005
R8250 a_22203_n358.n4 a_22203_n358.t7 3.6005
R8251 a_22203_n358.n3 a_22203_n358.t5 3.6005
R8252 a_22203_n358.n3 a_22203_n358.t6 3.6005
R8253 a_22203_n358.n0 a_22203_n358.n1 2.59067
R8254 a_22203_n358.n0 a_22203_n358.n8 2.22925
R8255 a_22203_n358.n2 a_22203_n358.t0 2.06607
R8256 a_22203_n358.n12 a_22203_n358.t2 2.06607
R8257 a_22203_n358.n2 a_22203_n358.t1 1.4923
R8258 a_22203_n358.t3 a_22203_n358.n12 1.4923
R8259 CLK.n0 CLK.t1 17.5205
R8260 CLK CLK.n0 13.2835
R8261 CLK.n0 CLK.t0 11.5588
R8262 a_n4208_n141.n2 a_n4208_n141.t4 26.5147
R8263 a_n4208_n141.n1 a_n4208_n141.t3 25.076
R8264 a_n4208_n141.n1 a_n4208_n141.t6 25.076
R8265 a_n4208_n141.n3 a_n4208_n141.t7 25.076
R8266 a_n4208_n141.n3 a_n4208_n141.t8 25.076
R8267 a_n4208_n141.n2 a_n4208_n141.t5 25.076
R8268 a_n4208_n141.n0 a_n4208_n141.t0 23.009
R8269 a_n4208_n141.n0 a_n4208_n141.t1 12.3005
R8270 a_n4208_n141.t2 a_n4208_n141.n1 11.2556
R8271 a_n4208_n141.n1 a_n4208_n141.n0 3.08843
R8272 a_n4208_n141.n1 a_n4208_n141.n3 2.8778
R8273 a_n4208_n141.n3 a_n4208_n141.n2 2.8778
R8274 a_n8471_219.n1 a_n8471_219.t6 31.1854
R8275 a_n8471_219.n0 a_n8471_219.t8 30.4809
R8276 a_n8471_219.n0 a_n8471_219.t7 29.7468
R8277 a_n8471_219.n0 a_n8471_219.t5 29.7468
R8278 a_n8471_219.n2 a_n8471_219.t10 29.7468
R8279 a_n8471_219.n2 a_n8471_219.t11 29.7468
R8280 a_n8471_219.n1 a_n8471_219.t9 29.7468
R8281 a_n8471_219.n3 a_n8471_219.t0 28.2414
R8282 a_n8471_219.n0 a_n8471_219.t3 11.7439
R8283 a_n8471_219.n3 a_n8471_219.t1 8.52921
R8284 a_n8471_219.n4 a_n8471_219.t4 4.50971
R8285 a_n8471_219.t2 a_n8471_219.n4 4.38259
R8286 a_n8471_219.n4 a_n8471_219.n0 3.32162
R8287 a_n8471_219.n0 a_n8471_219.n2 2.8778
R8288 a_n8471_219.n2 a_n8471_219.n1 2.8778
R8289 a_n8471_219.n0 a_n8471_219.n3 2.4541
R8290 a_23620_8319.n0 a_23620_8319.t5 56.5589
R8291 a_23620_8319.n1 a_23620_8319.t4 54.6195
R8292 a_23620_8319.n1 a_23620_8319.t3 54.3444
R8293 a_23620_8319.n0 a_23620_8319.t6 54.3444
R8294 a_23620_8319.n3 a_23620_8319.n2 7.32981
R8295 a_23620_8319.n3 a_23620_8319.n1 3.5139
R8296 a_23620_8319.t1 a_23620_8319.n3 1.76266
R8297 a_23620_8319.n2 a_23620_8319.t0 1.6385
R8298 a_23620_8319.n2 a_23620_8319.t2 1.6385
R8299 a_23620_8319.n1 a_23620_8319.n0 1.3316
R8300 a_n8537_n1530.n2 a_n8537_n1530.t13 48.7058
R8301 a_n8537_n1530.n10 a_n8537_n1530.t14 47.5611
R8302 a_n8537_n1530.t6 a_n8537_n1530.n11 47.5611
R8303 a_n8537_n1530.n7 a_n8537_n1530.t5 46.602
R8304 a_n8537_n1530.n6 a_n8537_n1530.t9 46.602
R8305 a_n8537_n1530.n5 a_n8537_n1530.t7 46.602
R8306 a_n8537_n1530.n4 a_n8537_n1530.t12 46.602
R8307 a_n8537_n1530.n3 a_n8537_n1530.t10 46.602
R8308 a_n8537_n1530.n2 a_n8537_n1530.t15 46.602
R8309 a_n8537_n1530.n0 a_n8537_n1530.n13 37.0921
R8310 a_n8537_n1530.t14 a_n8537_n1530.n9 33.9289
R8311 a_n8537_n1530.n12 a_n8537_n1530.t6 33.9289
R8312 a_n8537_n1530.n12 a_n8537_n1530.t11 28.7581
R8313 a_n8537_n1530.n11 a_n8537_n1530.t11 28.7581
R8314 a_n8537_n1530.t4 a_n8537_n1530.n9 28.7581
R8315 a_n8537_n1530.n10 a_n8537_n1530.t4 28.7581
R8316 a_n8537_n1530.n11 a_n8537_n1530.n10 18.8035
R8317 a_n8537_n1530.n17 a_n8537_n1530.t0 6.3005
R8318 a_n8537_n1530.n17 a_n8537_n1530.n16 4.85375
R8319 a_n8537_n1530.n15 a_n8537_n1530.n14 4.5005
R8320 a_n8537_n1530.n1 a_n8537_n1530.n0 1.83275
R8321 a_n8537_n1530.n13 a_n8537_n1530.n9 2.58592
R8322 a_n8537_n1530.n13 a_n8537_n1530.n12 2.58592
R8323 a_n8537_n1530.t3 a_n8537_n1530.n17 2.56843
R8324 a_n8537_n1530.t0 a_n8537_n1530.t1 1.6385
R8325 a_n8537_n1530.n16 a_n8537_n1530.n8 1.51412
R8326 a_n8537_n1530.n3 a_n8537_n1530.n2 1.00625
R8327 a_n8537_n1530.t2 a_n8537_n1530.t3 0.813
R8328 a_n8537_n1530.n7 a_n8537_n1530.n6 0.62375
R8329 a_n8537_n1530.n4 a_n8537_n1530.n3 0.57425
R8330 a_n8537_n1530.n6 a_n8537_n1530.n5 0.57425
R8331 a_n8537_n1530.n5 a_n8537_n1530.n4 0.25475
R8332 a_n8537_n1530.n14 a_n8537_n1530.n8 0.233801
R8333 a_n8537_n1530.n8 a_n8537_n1530.n7 0.169297
R8334 a_n8537_n1530.n15 a_n8537_n1530.n0 0.15575
R8335 a_n8537_n1530.n14 a_n8537_n1530.n1 0.148629
R8336 a_n8537_n1530.n16 a_n8537_n1530.n15 0.11975
R8337 a_n8537_n1530.n1 a_n8537_n1530.t8 46.6222
R8338 a_22115_253.n2 a_22115_253.t5 121.874
R8339 a_22115_253.t5 a_22115_253.t7 61.5152
R8340 a_22115_253.n0 a_22115_253.t4 52.378
R8341 a_22115_253.n0 a_22115_253.t3 17.7152
R8342 a_22115_253.n1 a_22115_253.t1 11.1158
R8343 a_22115_253.n1 a_22115_253.n2 9.95623
R8344 a_22115_253.n1 a_22115_253.n0 8.37615
R8345 a_22115_253.t0 a_22115_253.n1 8.02846
R8346 a_22115_253.n0 a_22115_253.t6 7.36133
R8347 a_22115_253.n2 a_22115_253.t2 6.7165
R8348 a_n8537_93.t4 a_n8537_93.n4 47.5611
R8349 a_n8537_93.n3 a_n8537_93.t12 47.5611
R8350 a_n8537_93.n0 a_n8537_93.n6 36.4925
R8351 a_n8537_93.n5 a_n8537_93.t4 33.9289
R8352 a_n8537_93.t12 a_n8537_93.n2 33.9289
R8353 a_n8537_93.n1 a_n8537_93.t3 31.0687
R8354 a_n8537_93.n0 a_n8537_93.t1 29.4084
R8355 a_n8537_93.n0 a_n8537_93.t14 29.3475
R8356 a_n8537_93.n0 a_n8537_93.t10 29.3475
R8357 a_n8537_93.n0 a_n8537_93.t5 29.3475
R8358 a_n8537_93.n0 a_n8537_93.t8 29.3475
R8359 a_n8537_93.n1 a_n8537_93.t6 29.3475
R8360 a_n8537_93.n1 a_n8537_93.t9 29.3475
R8361 a_n8537_93.n1 a_n8537_93.t7 29.3475
R8362 a_n8537_93.t11 a_n8537_93.n2 28.7581
R8363 a_n8537_93.n3 a_n8537_93.t11 28.7581
R8364 a_n8537_93.n5 a_n8537_93.t13 28.7581
R8365 a_n8537_93.n4 a_n8537_93.t13 28.7581
R8366 a_n8537_93.n4 a_n8537_93.n3 18.8035
R8367 a_n8537_93.n0 a_n8537_93.t2 10.616
R8368 a_n8537_93.t0 a_n8537_93.n0 4.49193
R8369 a_n8537_93.n0 a_n8537_93.n1 3.41375
R8370 a_n8537_93.n6 a_n8537_93.n2 2.58592
R8371 a_n8537_93.n6 a_n8537_93.n5 2.58592
R8372 CSVB.n10 CSVB.t21 50.888
R8373 CSVB.n11 CSVB.t19 50.888
R8374 CSVB.n12 CSVB.t29 50.888
R8375 CSVB.n13 CSVB.t23 50.888
R8376 CSVB.n14 CSVB.t18 50.888
R8377 CSVB.n15 CSVB.t24 50.888
R8378 CSVB.n16 CSVB.t20 50.888
R8379 CSVB.n17 CSVB.t22 50.888
R8380 CSVB.n10 CSVB.t4 50.888
R8381 CSVB.n11 CSVB.t8 50.888
R8382 CSVB.n12 CSVB.t12 50.888
R8383 CSVB.n13 CSVB.t0 50.888
R8384 CSVB.n14 CSVB.t10 50.888
R8385 CSVB.n15 CSVB.t14 50.888
R8386 CSVB.n16 CSVB.t6 50.888
R8387 CSVB.n17 CSVB.t2 50.888
R8388 CSVB.n44 CSVB.t25 29.0305
R8389 CSVB.n43 CSVB.t27 29.0305
R8390 CSVB.n47 CSVB.t28 28.988
R8391 CSVB.n45 CSVB.t26 28.988
R8392 CSVB.n49 CSVB.n48 2.2505
R8393 CSVB.n46 CSVB.n42 2.2505
R8394 CSVB.n18 CSVB.n17 2.05375
R8395 CSVB.n19 CSVB.n9 1.93679
R8396 CSVB.n2 CSVB.n1 1.53767
R8397 CSVB.n38 CSVB.n37 1.51597
R8398 CSVB.n4 CSVB.n3 1.51597
R8399 CSVB.n25 CSVB.n24 1.51597
R8400 CSVB.n44 CSVB.n42 1.16575
R8401 CSVB.n49 CSVB.n43 1.16575
R8402 CSVB CSVB.n50 0.662406
R8403 CSVB.n22 CSVB.n21 0.643357
R8404 CSVB.n23 CSVB.n7 0.643357
R8405 CSVB.n27 CSVB.n26 0.643357
R8406 CSVB.n28 CSVB.n6 0.643357
R8407 CSVB.n30 CSVB.n29 0.643357
R8408 CSVB.n31 CSVB.n5 0.643357
R8409 CSVB.n33 CSVB.n32 0.643357
R8410 CSVB.n35 CSVB.n34 0.643357
R8411 CSVB.n36 CSVB.n0 0.643357
R8412 CSVB.n40 CSVB.n39 0.643357
R8413 CSVB.n20 CSVB.n8 0.643357
R8414 CSVB.n1 CSVB.t9 0.3255
R8415 CSVB.n1 CSVB.t5 0.3255
R8416 CSVB.n37 CSVB.t1 0.3255
R8417 CSVB.n37 CSVB.t13 0.3255
R8418 CSVB.n3 CSVB.t15 0.3255
R8419 CSVB.n3 CSVB.t11 0.3255
R8420 CSVB.n24 CSVB.t3 0.3255
R8421 CSVB.n24 CSVB.t7 0.3255
R8422 CSVB.n9 CSVB.t16 0.293
R8423 CSVB.n9 CSVB.t17 0.293
R8424 CSVB.n40 CSVB.n2 0.176326
R8425 CSVB CSVB.n41 0.109022
R8426 CSVB.n20 CSVB.n19 0.0780912
R8427 CSVB.n19 CSVB.n18 0.0595326
R8428 CSVB.n48 CSVB.n46 0.04025
R8429 CSVB.n45 CSVB.n44 0.039655
R8430 CSVB.n47 CSVB.n43 0.039655
R8431 CSVB.n17 CSVB.n16 0.0352143
R8432 CSVB.n16 CSVB.n15 0.0352143
R8433 CSVB.n15 CSVB.n14 0.0352143
R8434 CSVB.n14 CSVB.n13 0.0352143
R8435 CSVB.n12 CSVB.n11 0.0352143
R8436 CSVB.n11 CSVB.n10 0.0352143
R8437 CSVB.n13 CSVB.n12 0.0352143
R8438 CSVB.n38 CSVB.n2 0.021882
R8439 CSVB.n46 CSVB.n45 0.021125
R8440 CSVB.n48 CSVB.n47 0.021125
R8441 CSVB.n50 CSVB.n42 0.020375
R8442 CSVB.n50 CSVB.n49 0.020375
R8443 CSVB.n22 CSVB.n8 0.0120888
R8444 CSVB.n23 CSVB.n22 0.0120888
R8445 CSVB.n26 CSVB.n23 0.0120888
R8446 CSVB.n30 CSVB.n6 0.0120888
R8447 CSVB.n31 CSVB.n30 0.0120888
R8448 CSVB.n32 CSVB.n31 0.0120888
R8449 CSVB.n36 CSVB.n35 0.0120888
R8450 CSVB.n39 CSVB.n36 0.0120888
R8451 CSVB.n21 CSVB.n20 0.0120888
R8452 CSVB.n21 CSVB.n7 0.0120888
R8453 CSVB.n27 CSVB.n7 0.0120888
R8454 CSVB.n28 CSVB.n27 0.0120888
R8455 CSVB.n29 CSVB.n28 0.0120888
R8456 CSVB.n29 CSVB.n5 0.0120888
R8457 CSVB.n33 CSVB.n5 0.0120888
R8458 CSVB.n34 CSVB.n33 0.0120888
R8459 CSVB.n34 CSVB.n0 0.0120888
R8460 CSVB.n41 CSVB.n40 0.0119019
R8461 CSVB.n26 CSVB.n25 0.0093785
R8462 CSVB.n35 CSVB.n4 0.0093785
R8463 CSVB.n39 CSVB.n38 0.00816355
R8464 CSVB.n18 CSVB.n8 0.00433245
R8465 CSVB.n25 CSVB.n6 0.00321028
R8466 CSVB.n32 CSVB.n4 0.00321028
R8467 CSVB.n41 CSVB.n0 0.000686916
R8468 DOWN.n4 DOWN.t2 47.5611
R8469 DOWN.n5 DOWN.t5 36.5005
R8470 DOWN.n2 DOWN.t9 33.21
R8471 DOWN.n1 DOWN.t4 33.21
R8472 DOWN.n4 DOWN.t6 28.7581
R8473 DOWN.n6 DOWN.n4 26.2141
R8474 DOWN.n5 DOWN.t8 17.6975
R8475 DOWN.n2 DOWN.t3 17.6975
R8476 DOWN.n1 DOWN.t7 17.6975
R8477 DOWN.n6 DOWN.n5 10.7293
R8478 DOWN.n0 DOWN.t1 9.96025
R8479 DOWN DOWN.n0 8.34205
R8480 DOWN.n7 DOWN.n6 8.0005
R8481 DOWN.n3 DOWN.n1 7.75675
R8482 DOWN.n3 DOWN.n2 7.75675
R8483 DOWN.n0 DOWN.t0 4.28587
R8484 DOWN.n7 DOWN.n3 3.21483
R8485 DOWN DOWN.n7 2.55187
R8486 a_21506_13215.n2 a_21506_13215.t10 51.0134
R8487 a_21506_13215.n2 a_21506_13215.t11 50.7576
R8488 a_21506_13215.n0 a_21506_13215.n1 1.90384
R8489 a_21506_13215.n7 a_21506_13215.n5 1.55709
R8490 a_21506_13215.n7 a_21506_13215.n6 1.51597
R8491 a_21506_13215.n4 a_21506_13215.n3 1.51597
R8492 a_21506_13215.n9 a_21506_13215.n8 1.51457
R8493 a_21506_13215.n0 a_21506_13215.n2 2.67807
R8494 a_21506_13215.n5 a_21506_13215.t8 0.3255
R8495 a_21506_13215.n5 a_21506_13215.t6 0.3255
R8496 a_21506_13215.n6 a_21506_13215.t4 0.3255
R8497 a_21506_13215.n6 a_21506_13215.t2 0.3255
R8498 a_21506_13215.n3 a_21506_13215.t5 0.3255
R8499 a_21506_13215.n3 a_21506_13215.t7 0.3255
R8500 a_21506_13215.n9 a_21506_13215.t3 0.3255
R8501 a_21506_13215.t9 a_21506_13215.n9 0.3255
R8502 a_21506_13215.n1 a_21506_13215.t1 0.293
R8503 a_21506_13215.n1 a_21506_13215.t0 0.293
R8504 a_21506_13215.n8 a_21506_13215.n4 0.0406869
R8505 a_21506_13215.n8 a_21506_13215.n7 0.0402196
R8506 a_21506_13215.n4 a_21506_13215.n0 0.171403
R8507 UP.n3 UP.t7 47.5611
R8508 UP.n0 UP.t4 44.2706
R8509 UP.n1 UP.t8 44.2706
R8510 UP.n4 UP.t2 36.5005
R8511 UP.n3 UP.t5 28.7581
R8512 UP.n0 UP.t9 28.7581
R8513 UP.n1 UP.t3 28.7581
R8514 UP.n5 UP.n4 26.2141
R8515 UP.n4 UP.t6 17.6975
R8516 UP.n5 UP.n3 10.7293
R8517 UP.n7 UP.t0 9.96082
R8518 UP.n6 UP.n5 8.4865
R8519 UP.n2 UP.n0 7.75675
R8520 UP.n2 UP.n1 7.75675
R8521 UP UP.n7 4.85216
R8522 UP.n7 UP.t1 4.28533
R8523 UP.n6 UP.n2 2.72883
R8524 UP UP.n6 2.41659
R8525 a_22941_7733.n0 a_22941_7733.t5 42.2199
R8526 a_22941_7733.n1 a_22941_7733.t0 40.4081
R8527 a_22941_7733.n0 a_22941_7733.t6 40.4081
R8528 a_22941_7733.n0 a_22941_7733.t4 40.4081
R8529 a_22941_7733.n0 a_22941_7733.t3 40.4081
R8530 a_22941_7733.t2 a_22941_7733.n1 7.4853
R8531 a_22941_7733.n1 a_22941_7733.t1 5.40883
R8532 a_22941_7733.n1 a_22941_7733.n0 2.96695
R8533 a_22115_1610.n2 a_22115_1610.t7 121.874
R8534 a_22115_1610.t7 a_22115_1610.t4 61.5152
R8535 a_22115_1610.n0 a_22115_1610.t3 52.378
R8536 a_22115_1610.n0 a_22115_1610.t5 17.7882
R8537 a_22115_1610.n1 a_22115_1610.t1 11.1158
R8538 a_22115_1610.n1 a_22115_1610.n2 9.95623
R8539 a_22115_1610.n1 a_22115_1610.n0 8.37615
R8540 a_22115_1610.t0 a_22115_1610.n1 8.02846
R8541 a_22115_1610.n0 a_22115_1610.t2 7.3005
R8542 a_22115_1610.n2 a_22115_1610.t6 6.7165
R8543 a_22115_n302.n2 a_22115_n302.t7 121.874
R8544 a_22115_n302.t7 a_22115_n302.t4 61.5152
R8545 a_22115_n302.n0 a_22115_n302.t2 52.378
R8546 a_22115_n302.n0 a_22115_n302.t3 17.7882
R8547 a_22115_n302.n1 a_22115_n302.t1 11.1158
R8548 a_22115_n302.n1 a_22115_n302.n2 9.95623
R8549 a_22115_n302.n1 a_22115_n302.n0 8.37615
R8550 a_22115_n302.t0 a_22115_n302.n1 8.02846
R8551 a_22115_n302.n0 a_22115_n302.t6 7.3005
R8552 a_22115_n302.n2 a_22115_n302.t5 6.7165
R8553 a_22388_3950.t1 a_22388_3950.n1 21.2275
R8554 a_22388_3950.n1 a_22388_3950.t5 18.9805
R8555 a_22388_3950.n0 a_22388_3950.t4 17.5205
R8556 a_22388_3950.n0 a_22388_3950.t2 11.5588
R8557 a_22388_3950.n1 a_22388_3950.t3 11.4372
R8558 a_22388_3950.t1 a_22388_3950.t0 8.60523
R8559 a_22388_3950.t1 a_22388_3950.n0 8.27396
C0 a_5840_13333 OUT 0.021787f
C1 a_25265_7733 VDD 1.11074f
C2 a_22963_1518 a_25675_477 0.010299f
C3 a_10825_n1138 VDD 0.119269f
C4 a_23455_n345 a_23083_n301 0.107446f
C5 a_22527_n715 a_24383_n345 0.023074f
C6 a_22527_1197 VDD 1.11698f
C7 a_21855_n1258 VDD 1.02007f
C8 a_22115_4951 a_22563_4951 0.013276f
C9 a_23508_2038 a_25334_3994 0.010314f
C10 a_25095_7733 VDD 0.02907f
C11 a_22963_1518 a_24383_217 0.24646f
C12 a_25587_574 a_25675_n394 0.010569f
C13 a_6993_n1138 VDD 0.119269f
C14 a_22527_n715 a_23083_n301 0.839895f
C15 a_3149_2840 a_3345_2840 0.099479f
C16 VDD LF 1.91842f
C17 a_21755_1082 a_22948_2038 0.060492f
C18 a_27014_14933 a_27814_14933 0.017628f
C19 a_22963_1518 a_24090_629 0.051285f
C20 a_23691_7733 VDD 0.82092f
C21 a_3161_n1138 VDD 0.119269f
C22 a_22527_n715 a_23455_n345 1.16391f
C23 a_26115_6933 OUT 0.131726f
C24 a_21667_4951 a_22115_4951 0.013276f
C25 a_1712_10253 a_1712_9373 0.016713f
C26 a_24755_6933 VDD 1.07973f
C27 a_22963_1518 a_23083_261 0.045667f
C28 a_n671_n1138 VDD 0.119269f
C29 a_21855_1126 VDD 0.827537f
C30 a_25265_7733 OUT 1.35531f
C31 a_3149_2840 a_n487_2840 0.072091f
C32 a_26049_6873 UP 0.024796f
C33 a_21755_1082 a_21855_2486 0.517726f
C34 a_22864_2486 a_24655_2486 0.232395f
C35 a_22963_1518 a_23455_217 0.026991f
C36 a_5840_8933 OUT 0.021174f
C37 a_n8659_n1230 VDD 0.38527f
C38 a_25587_n302 VDD 0.361712f
C39 a_n683_2840 a_n487_2840 0.099479f
C40 a_24207_4398 a_24655_4398 0.480927f
C41 a_22864_2486 a_24207_2486 0.099075f
C42 a_25675_1518 a_25587_1610 0.285629f
C43 a_22963_1518 a_22963_217 0.154909f
C44 VDD CSVB 11.8692f
C45 a_18673_2840 VDD 0.347176f
C46 a_22963_217 a_23423_n1258 0.016718f
C47 a_23691_7733 OUT 0.156974f
C48 a_25675_n394 VDD 0.131342f
C49 a_26115_6933 UP 0.266123f
C50 a_23508_2038 a_24655_4398 0.05477f
C51 a_22304_2486 a_24207_2486 0.524f
C52 a_22864_2486 a_22948_2038 0.827579f
C53 a_22963_1518 a_22527_574 0.098711f
C54 a_11009_2840 VDD 0.629273f
C55 a_24755_6933 OUT 0.529591f
C56 a_25265_7733 UP 0.180056f
C57 a_22864_4398 a_24655_4398 0.224841f
C58 a_23508_2038 a_24207_4398 0.050704f
C59 a_1220_13333 a_1220_12453 0.041784f
C60 a_22304_2486 a_22948_2038 0.318976f
C61 a_n2908_10253 a_n2908_9373 0.016713f
C62 a_7177_2840 VDD 0.629273f
C63 a_22864_4398 a_24207_4398 0.097396f
C64 a_5840_14213 OUT 0.056192f
C65 a_18477_2840 VDD 0.298308f
C66 a_21667_n786 a_21755_n830 0.285629f
C67 OUT CSVB 0.1832f
C68 VDD DOWN 1.15299f
C69 a_22864_4398 a_23508_2038 1.28745f
C70 a_22304_4398 a_24655_4398 0.041108f
C71 a_22304_2486 a_21855_2486 0.051973f
C72 a_21855_1126 a_22963_217 0.147928f
C73 a_3345_2840 VDD 0.629273f
C74 a_24655_2486 VDD 0.443621f
C75 a_24090_n669 VDD 0.371422f
C76 a_24755_6933 UP 1.50376f
C77 a_22304_4398 a_24207_4398 0.524441f
C78 a_22948_3950 a_23508_2038 0.542819f
C79 a_22304_2486 a_21755_1082 0.029378f
C80 a_21855_1126 a_22527_574 0.075252f
C81 a_14645_2840 VDD 0.298285f
C82 a_22963_217 a_25587_n302 0.025816f
C83 a_24207_2486 VDD 0.57564f
C84 a_24383_n345 VDD 0.524797f
C85 a_22948_3950 a_22864_4398 0.827579f
C86 a_22304_4398 a_23508_2038 0.290117f
C87 a_1712_8493 a_1712_7613 0.016713f
C88 a_n487_2840 VDD 0.629273f
C89 a_22948_2038 VDD 0.472672f
C90 a_23083_n301 VDD 0.397859f
C91 VDD VCTRL 6.47944f
C92 OUT DOWN 0.310357f
C93 LF FREERUN 2.375f
C94 a_22304_4398 a_22864_4398 0.79492f
C95 a_10813_2840 VDD 0.298285f
C96 a_24383_217 a_24383_n345 0.01024f
C97 a_23455_n345 VDD 0.186107f
C98 a_26049_6873 a_25265_6933 0.111757f
C99 a_22304_4398 a_22948_3950 0.318865f
C100 a_21855_2486 VDD 0.465743f
C101 a_22527_n715 VDD 1.11099f
C102 a_22304_2486 a_22864_2486 0.77678f
C103 a_6981_2840 VDD 0.298285f
C104 a_21755_1082 VDD 1.49699f
C105 a_26115_6933 a_25265_6933 0.394051f
C106 LF EX 0.037658f
C107 VDD CLK 0.697841f
C108 UP DOWN 0.487462f
C109 a_24383_1567 a_24090_1243 0.493186f
C110 a_n2908_8493 a_n2908_7613 0.016713f
C111 a_22963_217 a_24090_n669 0.05056f
C112 a_21755_n830 VDD 0.377188f
C113 a_25265_7733 a_25265_6933 0.09437f
C114 a_21855_4398 a_22304_4398 0.051973f
C115 a_23423_n1258 F6 1.62795f
C116 a_23795_3522 a_22304_2486 0.019418f
C117 a_5840_10693 a_5840_9813 0.016713f
C118 a_22963_217 a_24383_n345 0.266557f
C119 a_3149_2840 VDD 0.298285f
C120 a_21667_n786 VDD 0.278953f
C121 a_23347_3522 a_22304_2486 0.011215f
C122 a_23455_1567 a_24090_1243 0.021118f
C123 a_5840_8933 a_5840_8053 0.016713f
C124 a_n683_2840 VDD 0.298285f
C125 a_22963_217 a_23083_n301 0.032472f
C126 a_24891_4907 a_25339_4907 0.013103f
C127 a_23347_3522 a_23795_3522 0.012552f
C128 a_n9701_6193 VCTRL 0.073173f
C129 a_22963_1518 a_24090_1243 0.011266f
C130 a_22963_217 a_23455_n345 0.046461f
C131 a_22864_2486 VDD 1.09154f
C132 a_22527_1197 a_24090_1243 0.416346f
C133 a_22963_1518 a_24383_1567 0.014406f
C134 a_23455_1567 a_23083_1611 0.107446f
C135 a_22963_217 a_22527_n715 0.093423f
C136 a_22304_2486 VDD 1.48563f
C137 a_25587_574 VDD 0.222895f
C138 a_26115_6933 a_26049_6873 0.247434f
C139 a_23691_7733 a_23691_6933 0.022218f
C140 a_24443_4907 a_24891_4907 0.013103f
C141 a_1712_13773 a_1220_13333 0.016789f
C142 a_22899_3522 a_23347_3522 0.012552f
C143 a_23508_2038 a_25334_2082 0.010209f
C144 a_1220_10693 a_1220_9813 0.016713f
C145 a_22527_1197 a_24383_1567 0.023074f
C146 a_22963_1518 a_23083_1611 0.240887f
C147 a_25339_4907 VDD 0.337435f
C148 a_25675_477 a_25587_574 0.285629f
C149 a_24866_11400 CSVB 1.05249f
C150 a_23795_3522 VDD 0.340986f
C151 a_1220_13773 a_1220_13333 0.016789f
C152 a_22963_1518 a_23455_1567 0.018863f
C153 a_22527_1197 a_23083_1611 0.839895f
C154 a_1220_8933 a_1220_8053 0.016713f
C155 a_24891_4907 VDD 0.333625f
C156 a_23347_3522 VDD 0.332254f
C157 a_25265_7733 a_26795_7733 0.019086f
C158 FREERUN VCTRL 2.62362f
C159 a_23995_4907 a_24443_4907 0.013103f
C160 a_23883_3430 a_22304_2486 0.026153f
C161 a_22451_3522 a_22899_3522 0.012552f
C162 a_22527_1197 a_23455_1567 1.16391f
C163 a_24443_4907 VDD 0.331821f
C164 a_22899_3522 VDD 0.336412f
C165 a_25265_7733 a_26115_6933 1.15373f
C166 a_23883_3430 a_23795_3522 0.285629f
C167 a_22527_1197 a_22963_1518 0.280621f
C168 a_23995_4907 VDD 0.33177f
C169 a_22451_3522 VDD 0.343186f
C170 a_23547_4907 a_23995_4907 0.013103f
C171 a_25265_6933 DOWN 0.110426f
C172 a_23435_3430 a_23795_3522 0.086905f
C173 a_22003_3522 a_22451_3522 0.012222f
C174 a_23508_2038 DOWN 0.100842f
C175 a_23547_4907 VDD 0.332636f
C176 a_21667_574 a_21667_n786 0.010569f
C177 a_22003_3522 VDD 0.346078f
C178 a_25675_477 VDD 0.336735f
C179 a_21891_6933 CSVB 0.012207f
C180 a_25095_7733 a_25265_7733 0.019086f
C181 a_5840_14213 a_5840_13333 0.016713f
C182 VCTRL EX 14.052299f
C183 a_23435_3430 a_23347_3522 0.285629f
C184 a_23508_2038 a_24655_2486 0.057075f
C185 a_23099_4907 VDD 0.338717f
C186 a_21555_3522 VDD 0.404801f
C187 a_24383_217 VDD 0.520925f
C188 a_23099_4907 a_23547_4907 0.013103f
C189 a_25251_4951 a_25339_4907 0.285629f
C190 a_22987_3430 a_23347_3522 0.086905f
C191 a_21555_3522 a_22003_3522 0.012222f
C192 a_23508_2038 a_24207_2486 0.051499f
C193 a_1712_11133 a_1712_10253 0.016713f
C194 a_21855_1126 a_22963_1518 0.107397f
C195 a_22651_4907 VDD 0.337108f
C196 a_23883_3430 VDD 0.232629f
C197 a_24090_629 VDD 0.370377f
C198 a_24755_6933 a_25265_7733 0.183758f
C199 a_25251_4951 a_24891_4907 0.087174f
C200 a_25339_4907 UP 0.015573f
C201 a_18673_2840 a_18489_n1138 0.063905f
C202 a_23508_2038 a_22948_2038 0.542819f
C203 a_22987_3430 a_22899_3522 0.285629f
C204 VDD OUT 5.027411f
C205 a_24866_11400 a_27414_10401 0.023394f
C206 a_21855_1126 a_22527_1197 0.071077f
C207 a_1712_9373 a_1712_8493 0.016713f
C208 a_5840_10693 OUT 0.021174f
C209 a_22203_4907 VDD 0.342721f
C210 a_23435_3430 VDD 0.205239f
C211 a_23083_261 VDD 0.397896f
C212 a_24755_6933 a_25095_7733 0.012025f
C213 a_22651_4907 a_23099_4907 0.013103f
C214 a_24803_4951 a_24891_4907 0.285629f
C215 a_1220_13773 a_1712_13773 0.01254f
C216 a_22539_3430 a_22899_3522 0.086905f
C217 a_21755_1082 a_25587_1610 0.026006f
C218 a_21755_4907 VDD 0.396412f
C219 a_24090_629 a_24383_217 0.493186f
C220 a_22987_3430 VDD 0.208767f
C221 a_23455_217 VDD 0.186132f
C222 a_24803_4951 a_24443_4907 0.087174f
C223 a_11009_2840 a_14657_n1138 0.058694f
C224 a_26049_6873 DOWN 1.46893f
C225 a_22539_3430 a_22451_3522 0.285629f
C226 a_25251_4951 VDD 0.203335f
C227 a_22539_3430 VDD 0.212862f
C228 a_22963_217 VDD 0.58464f
C229 a_22203_4907 a_22651_4907 0.013103f
C230 a_24355_4951 a_24443_4907 0.285629f
C231 a_11009_2840 a_10825_n1138 0.046681f
C232 a_n9701_6193 VDD 0.588689f
C233 a_23508_2038 a_21755_1082 0.235746f
C234 a_23435_3430 a_23883_3430 0.013276f
C235 a_22091_3430 a_22451_3522 0.086742f
C236 a_n2908_11133 a_n2908_10253 0.016713f
C237 a_24803_4951 VDD 0.203482f
C238 VDD UP 1.20823f
C239 a_22091_3430 VDD 0.215751f
C240 a_22527_574 VDD 1.1139f
C241 a_24355_4951 a_23995_4907 0.087174f
C242 a_7177_2840 a_10825_n1138 0.058694f
C243 a_n2908_14213 a_n2908_13333 0.016713f
C244 a_26115_6933 DOWN 0.112163f
C245 a_22091_3430 a_22003_3522 0.285629f
C246 a_24355_4951 VDD 0.203482f
C247 a_n2908_9373 a_n2908_8493 0.016713f
C248 a_23455_217 a_24090_629 0.021118f
C249 a_22963_217 a_24383_217 0.015243f
C250 a_21643_3430 VDD 0.255715f
C251 a_21667_574 VDD 0.278953f
C252 a_21755_4907 a_22203_4907 0.013103f
C253 a_23907_4951 a_23995_4907 0.285629f
C254 a_7177_2840 a_6993_n1138 0.046681f
C255 a_25265_7733 DOWN 0.022257f
C256 a_22987_3430 a_23435_3430 0.013276f
C257 a_21643_3430 a_22003_3522 0.086742f
C258 a_5840_11573 a_5840_10693 0.016713f
C259 a_23907_4951 VDD 0.203482f
C260 a_22527_574 a_24383_217 0.023074f
C261 a_23455_217 a_23083_261 0.107446f
C262 a_22963_217 a_24090_629 0.010957f
C263 a_23907_4951 a_23547_4907 0.087174f
C264 a_n2908_14213 LF 0.030954f
C265 a_21643_3430 a_21555_3522 0.285629f
C266 a_21755_1082 a_24090_1243 0.042898f
C267 a_23459_4951 VDD 0.203629f
C268 a_22963_217 a_23083_261 0.242122f
C269 a_22527_574 a_24090_629 0.416346f
C270 a_25675_n394 a_25587_n302 0.285629f
C271 a_21755_477 VDD 0.377703f
C272 VDD FREERUN 9.8079f
C273 OUT UP 0.488677f
C274 a_23459_4951 a_23547_4907 0.285629f
C275 a_3345_2840 a_6993_n1138 0.058694f
C276 a_23508_2038 a_22864_2486 0.873597f
C277 a_22539_3430 a_22987_3430 0.013276f
C278 a_21755_1082 a_24383_1567 0.249206f
C279 a_22527_574 a_23083_261 0.839895f
C280 a_22963_217 a_23455_217 0.01975f
C281 a_23011_4951 VDD 0.205777f
C282 a_23459_4951 a_23099_4907 0.087174f
C283 a_3345_2840 a_3161_n1138 0.046681f
C284 a_1712_14653 a_1712_13773 0.016713f
C285 a_24755_6933 DOWN 0.022154f
C286 a_22864_4398 a_22864_2486 0.013905f
C287 a_23508_2038 a_22304_2486 0.132024f
C288 a_21755_1082 a_23083_1611 0.025834f
C289 a_5840_11573 OUT 0.021174f
C290 a_22563_4951 VDD 0.208263f
C291 a_22527_574 a_23455_217 1.16391f
C292 a_21855_4398 CLK 0.4864f
C293 a_24803_4951 a_25251_4951 0.013276f
C294 a_23011_4951 a_23099_4907 0.285629f
C295 a_25251_4951 UP 0.012056f
C296 a_22091_3430 a_22539_3430 0.013276f
C297 a_1220_11573 a_1220_10693 0.016713f
C298 a_21755_1082 a_23455_1567 0.032377f
C299 a_22115_4951 VDD 0.219078f
C300 a_22527_574 a_22963_217 0.307596f
C301 a_23011_4951 a_22651_4907 0.087174f
C302 a_18477_2840 a_18673_2840 0.106065f
C303 a_n487_2840 a_3161_n1138 0.058694f
C304 a_7177_2840 a_11009_2840 0.971124f
C305 a_1220_14653 a_1220_13773 0.016713f
C306 VDD EX 1.373f
C307 LF VCTRL 14.5504f
C308 a_22304_4398 a_22864_2486 0.173051f
C309 a_21755_1082 a_22963_1518 0.137044f
C310 a_21667_4951 VDD 0.339057f
C311 a_24655_4398 VDD 0.444754f
C312 a_25587_1610 VDD 0.355683f
C313 a_24355_4951 a_24803_4951 0.013276f
C314 a_22563_4951 a_22651_4907 0.285629f
C315 a_n487_2840 a_n671_n1138 0.046681f
C316 a_22304_4398 a_22304_2486 0.01764f
C317 a_21643_3430 a_22091_3430 0.013276f
C318 a_21755_1082 a_22527_1197 0.090966f
C319 a_21855_1126 a_23083_n301 0.227561f
C320 a_25587_1610 a_25675_477 0.010569f
C321 a_24207_4398 VDD 0.573638f
C322 a_25675_1518 VDD 0.133852f
C323 a_22563_4951 a_22203_4907 0.087174f
C324 a_24866_11400 VDD 0.112967f
C325 a_23508_2038 VDD 1.7957f
C326 a_23907_4951 a_24355_4951 0.013276f
C327 a_22115_4951 a_22203_4907 0.285629f
C328 a_14645_2840 a_11009_2840 0.072091f
C329 a_3345_2840 a_7177_2840 0.971124f
C330 a_5840_9813 a_5840_8933 0.016713f
C331 a_21855_1126 a_22527_n715 0.421686f
C332 VDD F6 0.825656f
C333 a_22864_4398 VDD 1.01835f
C334 a_22115_4951 a_21755_4907 0.087174f
C335 a_1220_12453 a_1712_11133 0.016758f
C336 a_21755_1082 a_21855_1126 0.77448f
C337 a_21755_477 a_21667_574 0.285629f
C338 a_22948_3950 VDD 0.483755f
C339 a_21667_4951 a_21755_4907 0.285629f
C340 a_23459_4951 a_23907_4951 0.013276f
C341 a_23995_4907 a_22304_4398 0.011841f
C342 a_10813_2840 a_11009_2840 0.099479f
C343 a_22955_6933 VDD 0.017288f
C344 a_22963_1518 a_25587_574 0.023971f
C345 a_22304_4398 VDD 1.3581f
C346 a_24090_1243 VDD 0.372354f
C347 a_25265_6933 OUT 0.505363f
C348 a_10813_2840 a_7177_2840 0.072091f
C349 a_23508_2038 a_23435_3430 0.014853f
C350 a_22304_2486 a_22527_1197 0.010446f
C351 a_24207_2486 a_24655_2486 0.480927f
C352 a_5840_8053 OUT 0.021174f
C353 a_24383_n345 a_24090_n669 0.493186f
C354 a_24383_1567 VDD 0.523241f
C355 a_23011_4951 a_23459_4951 0.013276f
C356 a_n487_2840 a_3345_2840 0.971124f
C357 a_1220_14653 a_1712_14653 0.01254f
C358 a_1220_9813 a_1220_8933 0.016713f
C359 a_26049_6873 VDD 0.544082f
C360 a_21855_4398 VDD 0.466607f
C361 a_23083_1611 VDD 0.400846f
C362 a_23691_6933 OUT 0.140037f
C363 a_22651_4907 a_22304_4398 0.011676f
C364 a_6981_2840 a_7177_2840 0.099479f
C365 a_n2908_12013 a_n2908_11133 0.016713f
C366 a_26795_7733 VDD 0.02976f
C367 a_18489_n1138 VDD 0.119269f
C368 a_23455_n345 a_24090_n669 0.021118f
C369 a_23455_1567 VDD 0.186856f
C370 a_22955_6933 OUT 0.137981f
C371 a_22563_4951 a_23011_4951 0.013276f
C372 a_25265_6933 UP 0.090359f
C373 a_23508_2038 UP 0.011399f
C374 a_22948_3950 a_22987_3430 0.010389f
C375 a_1220_12453 a_1220_11573 0.024172f
C376 a_26115_6933 VDD 0.066159f
C377 a_14657_n1138 VDD 0.119269f
C378 a_22527_n715 a_24090_n669 0.416346f
C379 a_22963_1518 VDD 1.21408f
C380 a_21891_6933 OUT 0.137216f
C381 a_23423_n1258 VDD 1.92098f
C382 FREERUN EX 1.00652f
C383 a_25095_6933 UP 0.012946f
C384 a_6981_2840 a_3345_2840 0.072091f
C385 a_22864_4398 UP 0.013776f
C386 F6 VSS 0.956754f
C387 CLK VSS 0.542905f
C388 EX VSS 3.99463f
C389 VCTRL VSS 12.8205f
C390 FREERUN VSS 15.262243f
C391 DOWN VSS 4.36871f
C392 UP VSS 3.12935f
C393 CSVB VSS 9.49f
C394 OUT VSS 31.541714f
C395 LF VSS 49.024185f
C396 VDD VSS 0.355867p
C397 a_23423_n1258 VSS 2.97904f
C398 a_21855_n1258 VSS 1.5783f
C399 a_25587_n302 VSS 0.300869f
C400 a_25675_n394 VSS 0.553649f
C401 a_24090_n669 VSS 0.463372f
C402 a_24383_n345 VSS 0.847615f
C403 a_23083_n301 VSS 0.304138f
C404 a_23455_n345 VSS 0.42522f
C405 a_22527_n715 VSS 1.48041f
C406 a_21755_n830 VSS 0.253834f
C407 a_21667_n786 VSS 0.510899f
C408 a_25587_574 VSS 0.503354f
C409 a_25675_477 VSS 0.29293f
C410 a_24383_217 VSS 0.847727f
C411 a_24090_629 VSS 0.46342f
C412 a_23083_261 VSS 0.304138f
C413 a_23455_217 VSS 0.42522f
C414 a_22963_217 VSS 1.34533f
C415 a_22527_574 VSS 1.47988f
C416 a_21667_574 VSS 0.510899f
C417 a_21755_477 VSS 0.255908f
C418 a_25587_1610 VSS 0.300869f
C419 a_25675_1518 VSS 0.561365f
C420 a_24090_1243 VSS 0.468603f
C421 a_24383_1567 VSS 0.851182f
C422 a_23083_1611 VSS 0.30791f
C423 a_23455_1567 VSS 0.425059f
C424 a_22963_1518 VSS 0.669822f
C425 a_22527_1197 VSS 1.48233f
C426 a_21855_1126 VSS 0.731146f
C427 a_24655_2486 VSS 0.49929f
C428 a_24207_2486 VSS 0.52813f
C429 a_22948_2038 VSS 0.653228f
C430 a_21855_2486 VSS 0.487857f
C431 a_21755_1082 VSS 2.34133f
C432 a_22864_2486 VSS 1.32222f
C433 a_22304_2486 VSS 1.62693f
C434 a_23795_3522 VSS 0.291705f
C435 a_23347_3522 VSS 0.285378f
C436 a_22899_3522 VSS 0.286621f
C437 a_22451_3522 VSS 0.288647f
C438 a_22003_3522 VSS 0.288752f
C439 a_21555_3522 VSS 0.292965f
C440 a_23883_3430 VSS 0.496144f
C441 a_23435_3430 VSS 0.476403f
C442 a_22987_3430 VSS 0.478057f
C443 a_22539_3430 VSS 0.482501f
C444 a_22091_3430 VSS 0.482791f
C445 a_21643_3430 VSS 0.49561f
C446 a_24655_4398 VSS 0.501653f
C447 a_24207_4398 VSS 0.525166f
C448 a_23508_2038 VSS 3.34568f
C449 a_22864_4398 VSS 1.37341f
C450 a_22948_3950 VSS 0.663054f
C451 a_22304_4398 VSS 1.79445f
C452 a_21855_4398 VSS 0.486507f
C453 a_18489_n1138 VSS 0.583015f
C454 a_14657_n1138 VSS 0.59026f
C455 a_10825_n1138 VSS 0.59026f
C456 a_6993_n1138 VSS 0.59026f
C457 a_3161_n1138 VSS 0.59026f
C458 a_n671_n1138 VSS 0.59026f
C459 a_n8659_n1230 VSS 2.04194f
C460 a_18673_2840 VSS 1.12107f
C461 a_11009_2840 VSS 3.50221f
C462 a_7177_2840 VSS 3.50221f
C463 a_18477_2840 VSS 0.393424f
C464 a_3345_2840 VSS 3.50221f
C465 a_14645_2840 VSS 0.393424f
C466 a_n487_2840 VSS 3.48363f
C467 a_10813_2840 VSS 0.393424f
C468 a_6981_2840 VSS 0.393424f
C469 a_3149_2840 VSS 0.393424f
C470 a_n683_2840 VSS 0.393424f
C471 a_25339_4907 VSS 0.44212f
C472 a_24891_4907 VSS 0.284703f
C473 a_24443_4907 VSS 0.284815f
C474 a_23995_4907 VSS 0.284088f
C475 a_23547_4907 VSS 0.284758f
C476 a_23099_4907 VSS 0.285892f
C477 a_22651_4907 VSS 0.283647f
C478 a_22203_4907 VSS 0.28405f
C479 a_21755_4907 VSS 0.294904f
C480 a_25251_4951 VSS 0.502807f
C481 a_24803_4951 VSS 0.487275f
C482 a_24355_4951 VSS 0.489361f
C483 a_23907_4951 VSS 0.486164f
C484 a_23459_4951 VSS 0.487236f
C485 a_23011_4951 VSS 0.486282f
C486 a_22563_4951 VSS 0.48952f
C487 a_22115_4951 VSS 0.486149f
C488 a_21667_4951 VSS 0.52688f
C489 a_26795_6933 VSS 0.012152f
C490 a_25265_6933 VSS 0.681068f
C491 a_23691_6933 VSS 0.682074f
C492 a_22955_6933 VSS 0.677414f
C493 a_21891_6933 VSS 0.606695f
C494 a_26049_6873 VSS 1.20759f
C495 a_26115_6933 VSS 0.175429f
C496 a_25265_7733 VSS 0.166494f
C497 a_23691_7733 VSS 0.055944f
C498 a_24755_6933 VSS 0.642077f
C499 a_n9701_6193 VSS 2.79685f
C500 a_16431_6193 VSS 0.790553f
C501 a_1712_7613 VSS 0.768303f
C502 a_n2908_7613 VSS 0.821503f
C503 a_5840_8053 VSS 0.667177f
C504 a_1220_8053 VSS 0.755702f
C505 a_1712_8493 VSS 0.738449f
C506 a_n2908_8493 VSS 0.80006f
C507 a_5840_8933 VSS 0.666596f
C508 a_1220_8933 VSS 0.73827f
C509 a_1712_9373 VSS 0.738245f
C510 a_n2908_9373 VSS 0.798803f
C511 a_27814_14933 VSS 0.674688f
C512 a_27414_10401 VSS 0.658975f
C513 a_27014_14933 VSS 0.669913f
C514 a_5840_9813 VSS 0.666585f
C515 a_1220_9813 VSS 0.738245f
C516 a_1712_10253 VSS 0.738245f
C517 a_n2908_10253 VSS 0.800006f
C518 a_5840_10693 VSS 0.666585f
C519 a_1220_10693 VSS 0.738245f
C520 a_1712_11133 VSS 0.741641f
C521 a_n2908_11133 VSS 0.798351f
C522 a_5840_11573 VSS 0.677754f
C523 a_1220_11573 VSS 0.755665f
C524 a_1220_12453 VSS 0.933081f
C525 a_n2908_12013 VSS 0.809581f
C526 a_24866_11400 VSS 3.02217f
C527 a_1220_13333 VSS 0.921533f
C528 a_5840_13333 VSS 0.677754f
C529 a_n2908_13333 VSS 0.808528f
C530 a_1712_13773 VSS 0.741641f
C531 a_1220_13773 VSS 0.741701f
C532 a_5840_14213 VSS 0.666585f
C533 a_n2908_14213 VSS 0.799661f
C534 a_1712_14653 VSS 0.75376f
C535 a_1220_14653 VSS 0.755212f
C536 a_22388_3950.t1 VSS 1.25053f
C537 a_22388_3950.t0 VSS 0.048467f
C538 a_22388_3950.t4 VSS 0.077986f
C539 a_22388_3950.t2 VSS 0.042413f
C540 a_22388_3950.n0 VSS 0.079885f
C541 a_22388_3950.t5 VSS 0.078379f
C542 a_22388_3950.t3 VSS 0.060967f
C543 a_22388_3950.n1 VSS 0.46137f
C544 a_22115_n302.t6 VSS 0.043151f
C545 a_22115_n302.n0 VSS 0.221428f
C546 a_22115_n302.n1 VSS 0.803219f
C547 a_22115_n302.t2 VSS 0.144509f
C548 a_22115_n302.t3 VSS 0.127487f
C549 a_22115_n302.t1 VSS 0.047684f
C550 a_22115_n302.t5 VSS 0.020325f
C551 a_22115_n302.t4 VSS 0.127787f
C552 a_22115_n302.t7 VSS 0.401653f
C553 a_22115_n302.n2 VSS 0.257957f
C554 a_22115_n302.t0 VSS 0.1048f
C555 a_22115_1610.t2 VSS 0.041275f
C556 a_22115_1610.n0 VSS 0.211801f
C557 a_22115_1610.n1 VSS 0.768297f
C558 a_22115_1610.t3 VSS 0.138226f
C559 a_22115_1610.t5 VSS 0.121944f
C560 a_22115_1610.t1 VSS 0.045611f
C561 a_22115_1610.t6 VSS 0.019441f
C562 a_22115_1610.t4 VSS 0.122231f
C563 a_22115_1610.t7 VSS 0.38419f
C564 a_22115_1610.n2 VSS 0.246741f
C565 a_22115_1610.t0 VSS 0.100244f
C566 a_22941_7733.t2 VSS 0.178922f
C567 a_22941_7733.n0 VSS 1.87028f
C568 a_22941_7733.n1 VSS 0.91684f
C569 a_22941_7733.t5 VSS 0.157433f
C570 a_22941_7733.t3 VSS 0.137792f
C571 a_22941_7733.t4 VSS 0.137792f
C572 a_22941_7733.t6 VSS 0.137792f
C573 a_22941_7733.t0 VSS 0.036593f
C574 a_22941_7733.t1 VSS 0.026552f
C575 a_21506_13215.n0 VSS 1.78222f
C576 a_21506_13215.t3 VSS 0.036394f
C577 a_21506_13215.t1 VSS 0.036394f
C578 a_21506_13215.t0 VSS 0.036394f
C579 a_21506_13215.n1 VSS 0.113776f
C580 a_21506_13215.t10 VSS 0.124218f
C581 a_21506_13215.t11 VSS 0.123932f
C582 a_21506_13215.n2 VSS 0.219528f
C583 a_21506_13215.t5 VSS 0.036394f
C584 a_21506_13215.t7 VSS 0.036394f
C585 a_21506_13215.n3 VSS 0.12902f
C586 a_21506_13215.n4 VSS 1.39739f
C587 a_21506_13215.t8 VSS 0.036394f
C588 a_21506_13215.t6 VSS 0.036394f
C589 a_21506_13215.n5 VSS 0.1382f
C590 a_21506_13215.t4 VSS 0.036394f
C591 a_21506_13215.t2 VSS 0.036394f
C592 a_21506_13215.n6 VSS 0.12902f
C593 a_21506_13215.n7 VSS 0.897035f
C594 a_21506_13215.n8 VSS 0.55272f
C595 a_21506_13215.n9 VSS 0.129001f
C596 a_21506_13215.t9 VSS 0.036394f
C597 CSVB.n0 VSS 0.059807f
C598 CSVB.t9 VSS 0.028706f
C599 CSVB.t5 VSS 0.028706f
C600 CSVB.n1 VSS 0.104914f
C601 CSVB.n2 VSS 0.387725f
C602 CSVB.t15 VSS 0.028706f
C603 CSVB.t11 VSS 0.028706f
C604 CSVB.n3 VSS 0.101765f
C605 CSVB.n4 VSS 0.088973f
C606 CSVB.n5 VSS 0.117715f
C607 CSVB.n6 VSS 0.072622f
C608 CSVB.n7 VSS 0.117715f
C609 CSVB.n8 VSS 0.077815f
C610 CSVB.t16 VSS 0.028706f
C611 CSVB.t17 VSS 0.028706f
C612 CSVB.n9 VSS 0.12063f
C613 CSVB.t2 VSS 0.097898f
C614 CSVB.t6 VSS 0.097898f
C615 CSVB.t14 VSS 0.097898f
C616 CSVB.t10 VSS 0.097898f
C617 CSVB.t12 VSS 0.097898f
C618 CSVB.t8 VSS 0.097898f
C619 CSVB.t4 VSS 0.097898f
C620 CSVB.t21 VSS 0.097898f
C621 CSVB.n10 VSS 0.148897f
C622 CSVB.t19 VSS 0.097898f
C623 CSVB.n11 VSS 0.18754f
C624 CSVB.t29 VSS 0.097898f
C625 CSVB.n12 VSS 0.187569f
C626 CSVB.t0 VSS 0.097898f
C627 CSVB.t23 VSS 0.097898f
C628 CSVB.n13 VSS 0.199892f
C629 CSVB.t18 VSS 0.097898f
C630 CSVB.n14 VSS 0.18754f
C631 CSVB.t24 VSS 0.097898f
C632 CSVB.n15 VSS 0.18754f
C633 CSVB.t20 VSS 0.097898f
C634 CSVB.n16 VSS 0.18754f
C635 CSVB.t22 VSS 0.097898f
C636 CSVB.n17 VSS 0.264491f
C637 CSVB.n18 VSS 0.521504f
C638 CSVB.n19 VSS 2.21064f
C639 CSVB.n20 VSS 0.807685f
C640 CSVB.n21 VSS 0.117715f
C641 CSVB.n22 VSS 0.117715f
C642 CSVB.n23 VSS 0.117715f
C643 CSVB.t3 VSS 0.028706f
C644 CSVB.t7 VSS 0.028706f
C645 CSVB.n24 VSS 0.101765f
C646 CSVB.n25 VSS 0.088973f
C647 CSVB.n26 VSS 0.103949f
C648 CSVB.n27 VSS 0.117715f
C649 CSVB.n28 VSS 0.117715f
C650 CSVB.n29 VSS 0.117715f
C651 CSVB.n30 VSS 0.117715f
C652 CSVB.n31 VSS 0.117715f
C653 CSVB.n32 VSS 0.072622f
C654 CSVB.n33 VSS 0.117715f
C655 CSVB.n34 VSS 0.117715f
C656 CSVB.n35 VSS 0.103949f
C657 CSVB.n36 VSS 0.117715f
C658 CSVB.t1 VSS 0.028706f
C659 CSVB.t13 VSS 0.028706f
C660 CSVB.n37 VSS 0.101765f
C661 CSVB.n38 VSS 0.219211f
C662 CSVB.n39 VSS 0.097779f
C663 CSVB.n40 VSS 0.532364f
C664 CSVB.n41 VSS 0.370391f
C665 CSVB.n42 VSS 0.076714f
C666 CSVB.t27 VSS 0.042007f
C667 CSVB.n43 VSS 0.063068f
C668 CSVB.t25 VSS 0.042007f
C669 CSVB.n44 VSS 0.063068f
C670 CSVB.t26 VSS 0.041946f
C671 CSVB.n45 VSS 0.037947f
C672 CSVB.n46 VSS 0.019045f
C673 CSVB.t28 VSS 0.041946f
C674 CSVB.n47 VSS 0.037947f
C675 CSVB.n48 VSS 0.019045f
C676 CSVB.n49 VSS 0.076714f
C677 CSVB.n50 VSS 0.406664f
C678 a_n8537_93.n0 VSS 6.09595f
C679 a_n8537_93.n1 VSS 1.08916f
C680 a_n8537_93.t0 VSS 0.287725f
C681 a_n8537_93.t3 VSS 0.060225f
C682 a_n8537_93.t7 VSS 0.038171f
C683 a_n8537_93.t9 VSS 0.038171f
C684 a_n8537_93.t6 VSS 0.038171f
C685 a_n8537_93.t8 VSS 0.038171f
C686 a_n8537_93.t5 VSS 0.038171f
C687 a_n8537_93.t10 VSS 0.038171f
C688 a_n8537_93.t14 VSS 0.038171f
C689 a_n8537_93.t1 VSS 0.012232f
C690 a_n8537_93.n2 VSS 0.232035f
C691 a_n8537_93.t13 VSS 0.056513f
C692 a_n8537_93.t11 VSS 0.056513f
C693 a_n8537_93.t12 VSS 0.096345f
C694 a_n8537_93.n3 VSS 0.097801f
C695 a_n8537_93.n4 VSS 0.097801f
C696 a_n8537_93.t4 VSS 0.096345f
C697 a_n8537_93.n5 VSS 0.232035f
C698 a_n8537_93.n6 VSS 9.97896f
C699 a_n8537_93.t2 VSS 0.04316f
C700 a_22115_253.t6 VSS 0.042682f
C701 a_22115_253.n0 VSS 0.221505f
C702 a_22115_253.n1 VSS 0.803219f
C703 a_22115_253.t7 VSS 0.127787f
C704 a_22115_253.t5 VSS 0.401653f
C705 a_22115_253.t2 VSS 0.020325f
C706 a_22115_253.n2 VSS 0.257957f
C707 a_22115_253.t4 VSS 0.144509f
C708 a_22115_253.t3 VSS 0.127878f
C709 a_22115_253.t1 VSS 0.047684f
C710 a_22115_253.t0 VSS 0.1048f
C711 a_n8537_n1530.n0 VSS 4.12067f
C712 a_n8537_n1530.n1 VSS 0.157388f
C713 a_n8537_n1530.t3 VSS 0.165534f
C714 a_n8537_n1530.t13 VSS 0.057058f
C715 a_n8537_n1530.t15 VSS 0.043005f
C716 a_n8537_n1530.n2 VSS 0.627589f
C717 a_n8537_n1530.t10 VSS 0.043005f
C718 a_n8537_n1530.n3 VSS 0.17591f
C719 a_n8537_n1530.t12 VSS 0.043005f
C720 a_n8537_n1530.n4 VSS 0.106964f
C721 a_n8537_n1530.t7 VSS 0.043005f
C722 a_n8537_n1530.n5 VSS 0.106964f
C723 a_n8537_n1530.t9 VSS 0.043005f
C724 a_n8537_n1530.n6 VSS 0.140818f
C725 a_n8537_n1530.t5 VSS 0.043005f
C726 a_n8537_n1530.n7 VSS 0.110239f
C727 a_n8537_n1530.n8 VSS 0.030516f
C728 a_n8537_n1530.n9 VSS 0.1818f
C729 a_n8537_n1530.t11 VSS 0.044278f
C730 a_n8537_n1530.t4 VSS 0.044278f
C731 a_n8537_n1530.t14 VSS 0.075487f
C732 a_n8537_n1530.n10 VSS 0.076628f
C733 a_n8537_n1530.n11 VSS 0.076628f
C734 a_n8537_n1530.t6 VSS 0.075487f
C735 a_n8537_n1530.n12 VSS 0.1818f
C736 a_n8537_n1530.n13 VSS 9.222469f
C737 a_n8537_n1530.t8 VSS 0.043067f
C738 a_n8537_n1530.n14 VSS 0.0391f
C739 a_n8537_n1530.n15 VSS 0.021881f
C740 a_n8537_n1530.n16 VSS 0.150424f
C741 a_n8537_n1530.t0 VSS 0.040253f
C742 a_n8537_n1530.t1 VSS 0.013418f
C743 a_n8537_n1530.n17 VSS 0.225262f
C744 a_n8537_n1530.t2 VSS 0.030056f
C745 a_23620_8319.t1 VSS 0.230327f
C746 a_23620_8319.n0 VSS 1.12967f
C747 a_23620_8319.n1 VSS 0.948259f
C748 a_23620_8319.t0 VSS 0.02864f
C749 a_23620_8319.t2 VSS 0.02864f
C750 a_23620_8319.n2 VSS 0.085133f
C751 a_23620_8319.t5 VSS 0.160449f
C752 a_23620_8319.t6 VSS 0.141303f
C753 a_23620_8319.t3 VSS 0.141303f
C754 a_23620_8319.t4 VSS 0.142193f
C755 a_23620_8319.n3 VSS 0.564088f
C756 a_n8471_219.n0 VSS 4.02225f
C757 a_n8471_219.n1 VSS 1.52386f
C758 a_n8471_219.n2 VSS 1.96436f
C759 a_n8471_219.n3 VSS 0.450257f
C760 a_n8471_219.t4 VSS 0.052129f
C761 a_n8471_219.t2 VSS 0.050494f
C762 a_n8471_219.t1 VSS 0.017122f
C763 a_n8471_219.t0 VSS 0.010371f
C764 a_n8471_219.t8 VSS 0.016824f
C765 a_n8471_219.t6 VSS 0.040735f
C766 a_n8471_219.t9 VSS 0.014537f
C767 a_n8471_219.t11 VSS 0.014537f
C768 a_n8471_219.t10 VSS 0.014537f
C769 a_n8471_219.t5 VSS 0.014537f
C770 a_n8471_219.t7 VSS 0.014537f
C771 a_n8471_219.t3 VSS 0.031516f
C772 a_n8471_219.n4 VSS 0.6474f
C773 a_n4208_n141.n0 VSS 0.168853f
C774 a_n4208_n141.n1 VSS 2.09118f
C775 a_n4208_n141.n2 VSS 0.918953f
C776 a_n4208_n141.n3 VSS 1.17828f
C777 a_n4208_n141.t4 VSS 0.026767f
C778 a_n4208_n141.t2 VSS 0.069682f
C779 a_22203_n358.n0 VSS 0.603745f
C780 a_22203_n358.n1 VSS 1.31566f
C781 a_22203_n358.t2 VSS 0.018938f
C782 a_22203_n358.t0 VSS 0.018938f
C783 a_22203_n358.t1 VSS 0.013677f
C784 a_22203_n358.n2 VSS 0.032956f
C785 a_22203_n358.n3 VSS 0.010391f
C786 a_22203_n358.n4 VSS 0.014693f
C787 a_22203_n358.t15 VSS 0.054532f
C788 a_22203_n358.t18 VSS 0.035955f
C789 a_22203_n358.t11 VSS 0.020179f
C790 a_22203_n358.n5 VSS 0.096198f
C791 a_22203_n358.t17 VSS 0.035955f
C792 a_22203_n358.t10 VSS 0.020179f
C793 a_22203_n358.n6 VSS 0.062148f
C794 a_22203_n358.t14 VSS 0.035955f
C795 a_22203_n358.t13 VSS 0.020179f
C796 a_22203_n358.n7 VSS 0.065252f
C797 a_22203_n358.n8 VSS 0.041506f
C798 a_22203_n358.t12 VSS 0.025088f
C799 a_22203_n358.t9 VSS 0.026733f
C800 a_22203_n358.n9 VSS 0.058633f
C801 a_22203_n358.t8 VSS 0.026841f
C802 a_22203_n358.t16 VSS 0.024974f
C803 a_22203_n358.n10 VSS 0.048595f
C804 a_22203_n358.t20 VSS 0.025088f
C805 a_22203_n358.t19 VSS 0.026733f
C806 a_22203_n358.n11 VSS 0.048589f
C807 a_22203_n358.n12 VSS 0.037604f
C808 a_22203_n358.t3 VSS 0.013677f
C809 a_n17351_68.n0 VSS 9.0379f
C810 a_n17351_68.t1 VSS 0.054646f
C811 a_n17351_68.n1 VSS 0.03151f
C812 a_n17351_68.t25 VSS 0.021495f
C813 a_n17351_68.t10 VSS 0.021495f
C814 a_n17351_68.t26 VSS 0.021495f
C815 a_n17351_68.t22 VSS 0.021495f
C816 a_n17351_68.t29 VSS 0.021495f
C817 a_n17351_68.t24 VSS 0.021495f
C818 a_n17351_68.t31 VSS 0.021495f
C819 a_n17351_68.t18 VSS 0.021495f
C820 a_n17351_68.t33 VSS 0.021495f
C821 a_n17351_68.t2 VSS 0.021495f
C822 a_n17351_68.t28 VSS 0.021495f
C823 a_n17351_68.t38 VSS 0.021495f
C824 a_n17351_68.t20 VSS 0.021495f
C825 a_n17351_68.t32 VSS 0.021495f
C826 a_n17351_68.t13 VSS 0.021495f
C827 a_n17351_68.t30 VSS 0.021495f
C828 a_n17351_68.t23 VSS 0.021495f
C829 a_n17351_68.t36 VSS 0.021495f
C830 a_n17351_68.n2 VSS 0.038431f
C831 a_n17351_68.n3 VSS 0.038431f
C832 a_n17351_68.n4 VSS 0.038431f
C833 a_n17351_68.n5 VSS 0.038431f
C834 a_n17351_68.n6 VSS 0.038431f
C835 a_n17351_68.n7 VSS 0.038431f
C836 a_n17351_68.n8 VSS 0.038431f
C837 a_n17351_68.n9 VSS 0.054398f
C838 a_n17351_68.t35 VSS 0.049194f
C839 a_n17351_68.n10 VSS 0.046483f
C840 a_n17351_68.n11 VSS 0.033586f
C841 a_n17351_68.n12 VSS 0.033586f
C842 a_n17351_68.n13 VSS 0.033586f
C843 a_n17351_68.n14 VSS 0.033586f
C844 a_n17351_68.n15 VSS 0.033586f
C845 a_n17351_68.n16 VSS 0.033586f
C846 a_n17351_68.n17 VSS 0.033586f
C847 a_n17351_68.n18 VSS 0.033586f
C848 a_n17351_68.n19 VSS 0.033586f
C849 a_n17351_68.n20 VSS 0.033586f
C850 a_n17351_68.n21 VSS 0.033586f
C851 a_n17351_68.n22 VSS 0.033586f
C852 a_n17351_68.n23 VSS 0.033586f
C853 a_n17351_68.n24 VSS 0.033586f
C854 a_n17351_68.n25 VSS 0.033586f
C855 a_n17351_68.n26 VSS 0.033586f
C856 a_n17351_68.n27 VSS 0.046483f
C857 a_n17351_68.t27 VSS 0.049194f
C858 a_n17351_68.n28 VSS 0.054398f
C859 a_n17351_68.n29 VSS 0.038431f
C860 a_n17351_68.n30 VSS 0.038431f
C861 a_n17351_68.n31 VSS 0.038431f
C862 a_n17351_68.n32 VSS 0.038431f
C863 a_n17351_68.n33 VSS 0.038431f
C864 a_n17351_68.n34 VSS 0.038431f
C865 a_n17351_68.n35 VSS 0.038431f
C866 a_n17351_68.n36 VSS 0.03151f
C867 a_n17351_68.n37 VSS 0.573797f
C868 a_n17351_68.n38 VSS 0.044944f
C869 a_n17351_68.t5 VSS 0.048364f
C870 a_n17351_68.t4 VSS 0.048364f
C871 a_n17351_68.t41 VSS 0.048364f
C872 a_n17351_68.t19 VSS 0.048364f
C873 a_n17351_68.t17 VSS 0.048364f
C874 a_n17351_68.t16 VSS 0.048364f
C875 a_n17351_68.t11 VSS 0.048364f
C876 a_n17351_68.t7 VSS 0.048364f
C877 a_n17351_68.t6 VSS 0.048364f
C878 a_n17351_68.t9 VSS 0.048364f
C879 a_n17351_68.t14 VSS 0.048364f
C880 a_n17351_68.t15 VSS 0.048364f
C881 a_n17351_68.t37 VSS 0.048364f
C882 a_n17351_68.t39 VSS 0.048364f
C883 a_n17351_68.t40 VSS 0.048364f
C884 a_n17351_68.t3 VSS 0.048364f
C885 a_n17351_68.t8 VSS 0.048364f
C886 a_n17351_68.t12 VSS 0.048364f
C887 a_n17351_68.n39 VSS 0.051865f
C888 a_n17351_68.n40 VSS 0.051865f
C889 a_n17351_68.n41 VSS 0.051865f
C890 a_n17351_68.n42 VSS 0.051865f
C891 a_n17351_68.n43 VSS 0.051865f
C892 a_n17351_68.n44 VSS 0.051865f
C893 a_n17351_68.n45 VSS 0.051865f
C894 a_n17351_68.n46 VSS 0.083096f
C895 a_n17351_68.t34 VSS 0.073372f
C896 a_n17351_68.n47 VSS 0.074214f
C897 a_n17351_68.n48 VSS 0.047021f
C898 a_n17351_68.n49 VSS 0.047021f
C899 a_n17351_68.n50 VSS 0.047021f
C900 a_n17351_68.n51 VSS 0.047021f
C901 a_n17351_68.n52 VSS 0.047021f
C902 a_n17351_68.n53 VSS 0.047021f
C903 a_n17351_68.n54 VSS 0.047021f
C904 a_n17351_68.n55 VSS 0.047021f
C905 a_n17351_68.n56 VSS 0.047021f
C906 a_n17351_68.n57 VSS 0.047021f
C907 a_n17351_68.n58 VSS 0.047021f
C908 a_n17351_68.n59 VSS 0.047021f
C909 a_n17351_68.n60 VSS 0.047021f
C910 a_n17351_68.n61 VSS 0.047021f
C911 a_n17351_68.n62 VSS 0.047021f
C912 a_n17351_68.n63 VSS 0.047021f
C913 a_n17351_68.n64 VSS 0.074214f
C914 a_n17351_68.t21 VSS 0.073372f
C915 a_n17351_68.n65 VSS 0.083096f
C916 a_n17351_68.n66 VSS 0.051865f
C917 a_n17351_68.n67 VSS 0.051865f
C918 a_n17351_68.n68 VSS 0.051865f
C919 a_n17351_68.n69 VSS 0.051865f
C920 a_n17351_68.n70 VSS 0.051865f
C921 a_n17351_68.n71 VSS 0.051865f
C922 a_n17351_68.n72 VSS 0.051865f
C923 a_n17351_68.n73 VSS 0.044944f
C924 a_n17351_68.n74 VSS 0.235157f
C925 a_n17351_68.n75 VSS 0.644365f
C926 a_n17351_68.t0 VSS 0.228393f
C927 a_n558_2704.n0 VSS 0.695343f
C928 a_n558_2704.n1 VSS 0.092881f
C929 a_n558_2704.n2 VSS 1.047f
C930 a_n558_2704.t1 VSS 0.010311f
C931 a_n558_2704.n3 VSS 0.996038f
C932 a_n558_2704.t0 VSS 0.015962f
C933 LF.t0 VSS 0.012567f
C934 LF.t48 VSS 0.262536f
C935 LF.t49 VSS 0.262536f
C936 LF.t47 VSS 0.262536f
C937 LF.t41 VSS 0.262536f
C938 LF.t42 VSS 0.262536f
C939 LF.n2 VSS 1.64736f
C940 LF.n3 VSS 2.03442f
C941 LF.t43 VSS 0.262536f
C942 LF.t44 VSS 0.262536f
C943 LF.t50 VSS 0.262536f
C944 LF.t45 VSS 0.262536f
C945 LF.t46 VSS 0.262536f
C946 LF.n4 VSS 6.82482f
C947 LF.n5 VSS 2.93674f
C948 LF.n19 VSS 0.074193f
C949 LF.n23 VSS 0.025477f
C950 LF.n27 VSS 0.02554f
C951 LF.n30 VSS 0.02554f
C952 LF.n34 VSS 0.02554f
C953 LF.n39 VSS 0.02554f
C954 LF.n51 VSS 0.02554f
C955 LF.n58 VSS 0.02554f
C956 LF.n75 VSS 0.02554f
C957 LF.n97 VSS 0.02554f
C958 LF.n104 VSS 0.051111f
C959 LF.n109 VSS 0.011351f
C960 VCTRL.t80 VSS 0.16959f
C961 VCTRL.t66 VSS 0.427048f
C962 VCTRL.t8 VSS 0.112876f
C963 VCTRL.t41 VSS 0.066527f
C964 VCTRL.t73 VSS 0.066527f
C965 VCTRL.n0 VSS 0.324794f
C966 VCTRL.t7 VSS 0.022176f
C967 VCTRL.t17 VSS 0.022176f
C968 VCTRL.n1 VSS 0.064071f
C969 VCTRL.t56 VSS 0.066527f
C970 VCTRL.t45 VSS 0.066527f
C971 VCTRL.n2 VSS 0.324794f
C972 VCTRL.t4 VSS 0.022176f
C973 VCTRL.t14 VSS 0.022176f
C974 VCTRL.n3 VSS 0.064071f
C975 VCTRL.t44 VSS 0.066527f
C976 VCTRL.t63 VSS 0.066527f
C977 VCTRL.n4 VSS 0.324794f
C978 VCTRL.t11 VSS 0.022176f
C979 VCTRL.t18 VSS 0.022176f
C980 VCTRL.n5 VSS 0.064071f
C981 VCTRL.t74 VSS 0.066527f
C982 VCTRL.t43 VSS 0.066527f
C983 VCTRL.n6 VSS 0.324794f
C984 VCTRL.t12 VSS 0.022176f
C985 VCTRL.t6 VSS 0.022176f
C986 VCTRL.n7 VSS 0.064071f
C987 VCTRL.t77 VSS 0.066527f
C988 VCTRL.t58 VSS 0.066527f
C989 VCTRL.n8 VSS 0.324794f
C990 VCTRL.t16 VSS 0.022176f
C991 VCTRL.t3 VSS 0.022176f
C992 VCTRL.n9 VSS 0.064071f
C993 VCTRL.t57 VSS 0.066527f
C994 VCTRL.t46 VSS 0.066527f
C995 VCTRL.n10 VSS 0.324794f
C996 VCTRL.t0 VSS 0.022176f
C997 VCTRL.t9 VSS 0.022176f
C998 VCTRL.n11 VSS 0.064071f
C999 VCTRL.t69 VSS 0.066527f
C1000 VCTRL.t76 VSS 0.066527f
C1001 VCTRL.n12 VSS 0.324794f
C1002 VCTRL.t1 VSS 0.022176f
C1003 VCTRL.t10 VSS 0.022176f
C1004 VCTRL.n13 VSS 0.064071f
C1005 VCTRL.t75 VSS 0.066527f
C1006 VCTRL.t79 VSS 0.066527f
C1007 VCTRL.n14 VSS 0.324794f
C1008 VCTRL.t5 VSS 0.022176f
C1009 VCTRL.t15 VSS 0.022176f
C1010 VCTRL.n15 VSS 0.064071f
C1011 VCTRL.t72 VSS 0.066527f
C1012 VCTRL.t71 VSS 0.066527f
C1013 VCTRL.n16 VSS 0.324794f
C1014 VCTRL.t2 VSS 0.022176f
C1015 VCTRL.t19 VSS 0.022176f
C1016 VCTRL.n17 VSS 0.064071f
C1017 VCTRL.t59 VSS 0.427048f
C1018 VCTRL.t13 VSS 0.112876f
C1019 VCTRL.n18 VSS 0.927434f
C1020 VCTRL.n19 VSS 0.923262f
C1021 VCTRL.n20 VSS 0.909616f
C1022 VCTRL.n21 VSS 0.909616f
C1023 VCTRL.n22 VSS 0.909616f
C1024 VCTRL.n23 VSS 0.909616f
C1025 VCTRL.n24 VSS 0.909616f
C1026 VCTRL.n25 VSS 0.909616f
C1027 VCTRL.n26 VSS 0.909616f
C1028 VCTRL.n27 VSS 0.923262f
C1029 VCTRL.n28 VSS 2.61648f
C1030 VCTRL.t24 VSS 0.427048f
C1031 VCTRL.t67 VSS 0.112876f
C1032 VCTRL.t23 VSS 0.066527f
C1033 VCTRL.t35 VSS 0.066527f
C1034 VCTRL.n29 VSS 0.324794f
C1035 VCTRL.t62 VSS 0.022176f
C1036 VCTRL.t61 VSS 0.022176f
C1037 VCTRL.n30 VSS 0.064071f
C1038 VCTRL.t22 VSS 0.066527f
C1039 VCTRL.t28 VSS 0.066527f
C1040 VCTRL.n31 VSS 0.324794f
C1041 VCTRL.t50 VSS 0.022176f
C1042 VCTRL.t42 VSS 0.022176f
C1043 VCTRL.n32 VSS 0.064071f
C1044 VCTRL.t20 VSS 0.066527f
C1045 VCTRL.t26 VSS 0.066527f
C1046 VCTRL.n33 VSS 0.324794f
C1047 VCTRL.t52 VSS 0.022176f
C1048 VCTRL.t70 VSS 0.022176f
C1049 VCTRL.n34 VSS 0.064071f
C1050 VCTRL.t39 VSS 0.066527f
C1051 VCTRL.t32 VSS 0.066527f
C1052 VCTRL.n35 VSS 0.324794f
C1053 VCTRL.t64 VSS 0.022176f
C1054 VCTRL.t48 VSS 0.022176f
C1055 VCTRL.n36 VSS 0.064071f
C1056 VCTRL.t38 VSS 0.066527f
C1057 VCTRL.t30 VSS 0.066527f
C1058 VCTRL.n37 VSS 0.324794f
C1059 VCTRL.t40 VSS 0.022176f
C1060 VCTRL.t54 VSS 0.022176f
C1061 VCTRL.n38 VSS 0.064071f
C1062 VCTRL.t37 VSS 0.066527f
C1063 VCTRL.t29 VSS 0.066527f
C1064 VCTRL.n39 VSS 0.324794f
C1065 VCTRL.t78 VSS 0.022176f
C1066 VCTRL.t55 VSS 0.022176f
C1067 VCTRL.n40 VSS 0.064071f
C1068 VCTRL.t36 VSS 0.066527f
C1069 VCTRL.t31 VSS 0.066527f
C1070 VCTRL.n41 VSS 0.324794f
C1071 VCTRL.t60 VSS 0.022176f
C1072 VCTRL.t49 VSS 0.022176f
C1073 VCTRL.n42 VSS 0.064071f
C1074 VCTRL.t34 VSS 0.066527f
C1075 VCTRL.t21 VSS 0.066527f
C1076 VCTRL.n43 VSS 0.324794f
C1077 VCTRL.t53 VSS 0.022176f
C1078 VCTRL.t51 VSS 0.022176f
C1079 VCTRL.n44 VSS 0.064071f
C1080 VCTRL.t27 VSS 0.066527f
C1081 VCTRL.t25 VSS 0.066527f
C1082 VCTRL.n45 VSS 0.324794f
C1083 VCTRL.t68 VSS 0.022176f
C1084 VCTRL.t65 VSS 0.022176f
C1085 VCTRL.n46 VSS 0.064071f
C1086 VCTRL.t33 VSS 0.427048f
C1087 VCTRL.t47 VSS 0.112876f
C1088 VCTRL.n47 VSS 0.927434f
C1089 VCTRL.n48 VSS 0.923262f
C1090 VCTRL.n49 VSS 0.909616f
C1091 VCTRL.n50 VSS 0.909616f
C1092 VCTRL.n51 VSS 0.909616f
C1093 VCTRL.n52 VSS 0.909616f
C1094 VCTRL.n53 VSS 0.909616f
C1095 VCTRL.n54 VSS 0.909616f
C1096 VCTRL.n55 VSS 0.909616f
C1097 VCTRL.n56 VSS 0.923262f
C1098 VCTRL.n57 VSS 1.09418f
C1099 VCTRL.n58 VSS 2.24736f
C1100 EX.t32 VSS 0.054066f
C1101 EX.t28 VSS 0.054066f
C1102 EX.n0 VSS 0.248503f
C1103 EX.t17 VSS 0.018022f
C1104 EX.t3 VSS 0.018022f
C1105 EX.n1 VSS 0.081213f
C1106 EX.t39 VSS 0.054066f
C1107 EX.t33 VSS 0.054066f
C1108 EX.n2 VSS 0.248503f
C1109 EX.t13 VSS 0.018022f
C1110 EX.t6 VSS 0.018022f
C1111 EX.n3 VSS 0.081213f
C1112 EX.t37 VSS 0.054066f
C1113 EX.t36 VSS 0.054066f
C1114 EX.n4 VSS 0.248503f
C1115 EX.t18 VSS 0.018022f
C1116 EX.t5 VSS 0.018022f
C1117 EX.n5 VSS 0.081213f
C1118 EX.t24 VSS 0.054066f
C1119 EX.t31 VSS 0.054066f
C1120 EX.n6 VSS 0.248503f
C1121 EX.t11 VSS 0.018022f
C1122 EX.t15 VSS 0.018022f
C1123 EX.n7 VSS 0.081213f
C1124 EX.t27 VSS 0.054066f
C1125 EX.t26 VSS 0.054066f
C1126 EX.n8 VSS 0.248503f
C1127 EX.t7 VSS 0.018022f
C1128 EX.t14 VSS 0.018022f
C1129 EX.n9 VSS 0.081213f
C1130 EX.t21 VSS 0.054066f
C1131 EX.t38 VSS 0.054066f
C1132 EX.n10 VSS 0.248503f
C1133 EX.t8 VSS 0.018022f
C1134 EX.t0 VSS 0.018022f
C1135 EX.n11 VSS 0.081213f
C1136 EX.t29 VSS 0.054066f
C1137 EX.t35 VSS 0.054066f
C1138 EX.n12 VSS 0.248503f
C1139 EX.t16 VSS 0.018022f
C1140 EX.t2 VSS 0.018022f
C1141 EX.n13 VSS 0.081213f
C1142 EX.t23 VSS 0.054066f
C1143 EX.t22 VSS 0.054066f
C1144 EX.n14 VSS 0.248503f
C1145 EX.t12 VSS 0.018022f
C1146 EX.t19 VSS 0.018022f
C1147 EX.n15 VSS 0.081213f
C1148 EX.t34 VSS 0.054066f
C1149 EX.t25 VSS 0.054066f
C1150 EX.n16 VSS 0.248503f
C1151 EX.t1 VSS 0.018022f
C1152 EX.t4 VSS 0.018022f
C1153 EX.n17 VSS 0.081213f
C1154 EX.t30 VSS 0.054066f
C1155 EX.t20 VSS 0.054066f
C1156 EX.n18 VSS 0.248503f
C1157 EX.t10 VSS 0.018022f
C1158 EX.t9 VSS 0.018022f
C1159 EX.n19 VSS 0.081213f
C1160 EX.n20 VSS 0.791815f
C1161 EX.n21 VSS 0.881926f
C1162 EX.n22 VSS 0.881926f
C1163 EX.n23 VSS 0.881926f
C1164 EX.n24 VSS 0.881926f
C1165 EX.n25 VSS 0.881926f
C1166 EX.n26 VSS 0.881926f
C1167 EX.n27 VSS 0.881926f
C1168 EX.n28 VSS 0.881926f
C1169 EX.n29 VSS 2.13169f
C1170 FREERUN.n0 VSS 0.07358f
C1171 FREERUN.t37 VSS 0.079178f
C1172 FREERUN.t23 VSS 0.079178f
C1173 FREERUN.t40 VSS 0.079178f
C1174 FREERUN.t30 VSS 0.079178f
C1175 FREERUN.t4 VSS 0.079178f
C1176 FREERUN.t34 VSS 0.079178f
C1177 FREERUN.t7 VSS 0.079178f
C1178 FREERUN.t25 VSS 0.079178f
C1179 FREERUN.t12 VSS 0.079178f
C1180 FREERUN.t18 VSS 0.079178f
C1181 FREERUN.t3 VSS 0.079178f
C1182 FREERUN.t15 VSS 0.079178f
C1183 FREERUN.t27 VSS 0.079178f
C1184 FREERUN.t9 VSS 0.079178f
C1185 FREERUN.t24 VSS 0.079178f
C1186 FREERUN.t5 VSS 0.079178f
C1187 FREERUN.t32 VSS 0.079178f
C1188 FREERUN.t14 VSS 0.079178f
C1189 FREERUN.n1 VSS 0.08491f
C1190 FREERUN.n2 VSS 0.08491f
C1191 FREERUN.n3 VSS 0.08491f
C1192 FREERUN.n4 VSS 0.08491f
C1193 FREERUN.n5 VSS 0.08491f
C1194 FREERUN.n6 VSS 0.08491f
C1195 FREERUN.n7 VSS 0.08491f
C1196 FREERUN.n8 VSS 0.136038f
C1197 FREERUN.t13 VSS 0.12012f
C1198 FREERUN.n9 VSS 0.121498f
C1199 FREERUN.n10 VSS 0.076979f
C1200 FREERUN.n11 VSS 0.076979f
C1201 FREERUN.n12 VSS 0.076979f
C1202 FREERUN.n13 VSS 0.076979f
C1203 FREERUN.n14 VSS 0.076979f
C1204 FREERUN.n15 VSS 0.076979f
C1205 FREERUN.n16 VSS 0.076979f
C1206 FREERUN.n17 VSS 0.076979f
C1207 FREERUN.n18 VSS 0.076979f
C1208 FREERUN.n19 VSS 0.076979f
C1209 FREERUN.n20 VSS 0.076979f
C1210 FREERUN.n21 VSS 0.076979f
C1211 FREERUN.n22 VSS 0.076979f
C1212 FREERUN.n23 VSS 0.076979f
C1213 FREERUN.n24 VSS 0.076979f
C1214 FREERUN.n25 VSS 0.076979f
C1215 FREERUN.n26 VSS 0.121498f
C1216 FREERUN.t1 VSS 0.12012f
C1217 FREERUN.n27 VSS 0.136038f
C1218 FREERUN.n28 VSS 0.08491f
C1219 FREERUN.n29 VSS 0.08491f
C1220 FREERUN.n30 VSS 0.08491f
C1221 FREERUN.n31 VSS 0.08491f
C1222 FREERUN.n32 VSS 0.08491f
C1223 FREERUN.n33 VSS 0.08491f
C1224 FREERUN.n34 VSS 0.08491f
C1225 FREERUN.n35 VSS 0.07358f
C1226 FREERUN.n36 VSS 2.10553f
C1227 FREERUN.t38 VSS 0.041918f
C1228 FREERUN.n37 VSS 1.04593f
C1229 FREERUN.n38 VSS 0.051586f
C1230 FREERUN.t33 VSS 0.03519f
C1231 FREERUN.t41 VSS 0.03519f
C1232 FREERUN.t21 VSS 0.03519f
C1233 FREERUN.t39 VSS 0.03519f
C1234 FREERUN.t20 VSS 0.03519f
C1235 FREERUN.t29 VSS 0.03519f
C1236 FREERUN.t10 VSS 0.03519f
C1237 FREERUN.t36 VSS 0.03519f
C1238 FREERUN.t0 VSS 0.03519f
C1239 FREERUN.t8 VSS 0.03519f
C1240 FREERUN.t28 VSS 0.03519f
C1241 FREERUN.t17 VSS 0.03519f
C1242 FREERUN.t2 VSS 0.03519f
C1243 FREERUN.t19 VSS 0.03519f
C1244 FREERUN.t11 VSS 0.03519f
C1245 FREERUN.t31 VSS 0.03519f
C1246 FREERUN.t6 VSS 0.03519f
C1247 FREERUN.t26 VSS 0.03519f
C1248 FREERUN.n39 VSS 0.062916f
C1249 FREERUN.n40 VSS 0.062916f
C1250 FREERUN.n41 VSS 0.062916f
C1251 FREERUN.n42 VSS 0.062916f
C1252 FREERUN.n43 VSS 0.062916f
C1253 FREERUN.n44 VSS 0.062916f
C1254 FREERUN.n45 VSS 0.062916f
C1255 FREERUN.n46 VSS 0.089056f
C1256 FREERUN.t22 VSS 0.080537f
C1257 FREERUN.n47 VSS 0.076099f
C1258 FREERUN.n48 VSS 0.054985f
C1259 FREERUN.n49 VSS 0.054985f
C1260 FREERUN.n50 VSS 0.054985f
C1261 FREERUN.n51 VSS 0.054985f
C1262 FREERUN.n52 VSS 0.054985f
C1263 FREERUN.n53 VSS 0.054985f
C1264 FREERUN.n54 VSS 0.054985f
C1265 FREERUN.n55 VSS 0.054985f
C1266 FREERUN.n56 VSS 0.054985f
C1267 FREERUN.n57 VSS 0.054985f
C1268 FREERUN.n58 VSS 0.054985f
C1269 FREERUN.n59 VSS 0.054985f
C1270 FREERUN.n60 VSS 0.054985f
C1271 FREERUN.n61 VSS 0.054985f
C1272 FREERUN.n62 VSS 0.054985f
C1273 FREERUN.n63 VSS 0.054985f
C1274 FREERUN.n64 VSS 0.076099f
C1275 FREERUN.t16 VSS 0.080537f
C1276 FREERUN.n65 VSS 0.089056f
C1277 FREERUN.n66 VSS 0.062916f
C1278 FREERUN.n67 VSS 0.062916f
C1279 FREERUN.n68 VSS 0.062916f
C1280 FREERUN.n69 VSS 0.062916f
C1281 FREERUN.n70 VSS 0.062916f
C1282 FREERUN.n71 VSS 0.062916f
C1283 FREERUN.n72 VSS 0.062916f
C1284 FREERUN.n73 VSS 0.051586f
C1285 FREERUN.n74 VSS 2.10446f
C1286 FREERUN.t35 VSS 0.094642f
C1287 FREERUN.n75 VSS 1.10052f
C1288 FREERUN.n76 VSS 0.364432f
C1289 a_22388_2038.t1 VSS 1.25053f
C1290 a_22388_2038.t0 VSS 0.048467f
C1291 a_22388_2038.t5 VSS 0.077986f
C1292 a_22388_2038.t3 VSS 0.042413f
C1293 a_22388_2038.n0 VSS 0.079885f
C1294 a_22388_2038.t2 VSS 0.078379f
C1295 a_22388_2038.t4 VSS 0.060967f
C1296 a_22388_2038.n1 VSS 0.46137f
C1297 a_5840_7613.t1 VSS 26.4671f
C1298 a_5840_7613.t0 VSS 0.032928f
C1299 OUT.n50 VSS 0.013451f
C1300 OUT.n53 VSS 0.010406f
C1301 OUT.n56 VSS 0.019079f
C1302 OUT.n61 VSS 0.013472f
C1303 OUT.n70 VSS 0.031984f
C1304 OUT.t13 VSS 0.967121f
C1305 OUT.t12 VSS 0.967121f
C1306 OUT.t9 VSS 0.967121f
C1307 OUT.t18 VSS 0.967121f
C1308 OUT.t20 VSS 0.967121f
C1309 OUT.t11 VSS 0.967121f
C1310 OUT.n168 VSS 3.9853f
C1311 OUT.t10 VSS 0.967121f
C1312 OUT.t15 VSS 0.967121f
C1313 OUT.n169 VSS 4.471779f
C1314 OUT.t14 VSS 0.967121f
C1315 OUT.t16 VSS 0.967121f
C1316 OUT.n170 VSS 4.471779f
C1317 OUT.t19 VSS 0.967121f
C1318 OUT.t17 VSS 0.967121f
C1319 OUT.n171 VSS 4.68256f
C1320 OUT.n172 VSS 0.602413f
C1321 OUT.n173 VSS 0.012868f
C1322 VDD.n0 VSS 7.67727f
C1323 VDD.n2 VSS 0.070629f
C1324 VDD.n4 VSS 0.043242f
C1325 VDD.n5 VSS 0.066401f
C1326 VDD.n6 VSS 0.078621f
C1327 VDD.n7 VSS 0.078621f
C1328 VDD.n8 VSS 0.070165f
C1329 VDD.n9 VSS 0.04418f
C1330 VDD.n12 VSS 0.022784f
C1331 VDD.t168 VSS 0.02234f
C1332 VDD.n13 VSS 0.077567f
C1333 VDD.n14 VSS 0.298952f
C1334 VDD.n15 VSS 0.298952f
C1335 VDD.n16 VSS 0.025672f
C1336 VDD.n17 VSS 0.027158f
C1337 VDD.t167 VSS 0.200086f
C1338 VDD.n20 VSS 0.027158f
C1339 VDD.n21 VSS 0.015767f
C1340 VDD.n22 VSS 0.030221f
C1341 VDD.n23 VSS 0.051316f
C1342 VDD.n24 VSS 0.034539f
C1343 VDD.n29 VSS 0.018534f
C1344 VDD.n32 VSS 0.354208f
C1345 VDD.t216 VSS 0.159289f
C1346 VDD.t241 VSS 0.11513f
C1347 VDD.t242 VSS 0.11513f
C1348 VDD.t316 VSS 0.11513f
C1349 VDD.t270 VSS 0.11513f
C1350 VDD.t271 VSS 0.11513f
C1351 VDD.t240 VSS 0.11513f
C1352 VDD.t180 VSS 0.11513f
C1353 VDD.t213 VSS 0.11513f
C1354 VDD.t214 VSS 0.086347f
C1355 VDD.n33 VSS 0.057565f
C1356 VDD.t315 VSS 0.086347f
C1357 VDD.t177 VSS 0.11513f
C1358 VDD.t269 VSS 0.11513f
C1359 VDD.t217 VSS 0.11513f
C1360 VDD.t178 VSS 0.11513f
C1361 VDD.t179 VSS 0.11513f
C1362 VDD.t212 VSS 0.11513f
C1363 VDD.t243 VSS 0.11513f
C1364 VDD.t176 VSS 0.11513f
C1365 VDD.t239 VSS 0.159289f
C1366 VDD.n34 VSS 0.354208f
C1367 VDD.n35 VSS 0.011454f
C1368 VDD.n36 VSS 0.043242f
C1369 VDD.n37 VSS 0.112603f
C1370 VDD.n38 VSS 0.097652f
C1371 VDD.n39 VSS 0.043242f
C1372 VDD.n40 VSS 0.078621f
C1373 VDD.n41 VSS 0.078621f
C1374 VDD.n42 VSS 0.074393f
C1375 VDD.n43 VSS 0.080066f
C1376 VDD.n44 VSS 0.354208f
C1377 VDD.t157 VSS 0.159289f
C1378 VDD.t159 VSS 0.11513f
C1379 VDD.t201 VSS 0.11513f
C1380 VDD.t162 VSS 0.11513f
C1381 VDD.t166 VSS 0.11513f
C1382 VDD.t141 VSS 0.11513f
C1383 VDD.t161 VSS 0.11513f
C1384 VDD.t196 VSS 0.11513f
C1385 VDD.t312 VSS 0.11513f
C1386 VDD.t175 VSS 0.086347f
C1387 VDD.n45 VSS 0.057565f
C1388 VDD.t160 VSS 0.086347f
C1389 VDD.t158 VSS 0.11513f
C1390 VDD.t195 VSS 0.11513f
C1391 VDD.t202 VSS 0.11513f
C1392 VDD.t163 VSS 0.11513f
C1393 VDD.t313 VSS 0.11513f
C1394 VDD.t142 VSS 0.11513f
C1395 VDD.t299 VSS 0.11513f
C1396 VDD.t194 VSS 0.11513f
C1397 VDD.t193 VSS 0.159289f
C1398 VDD.n46 VSS 0.354208f
C1399 VDD.n54 VSS 0.034539f
C1400 VDD.n55 VSS 0.193776f
C1401 VDD.n56 VSS 2.27778f
C1402 VDD.n57 VSS 0.057934f
C1403 VDD.n58 VSS 0.018993f
C1404 VDD.t164 VSS 0.064126f
C1405 VDD.t91 VSS 0.099064f
C1406 VDD.t23 VSS 0.099064f
C1407 VDD.t39 VSS 0.099064f
C1408 VDD.t247 VSS 0.105034f
C1409 VDD.t255 VSS 0.064789f
C1410 VDD.t292 VSS 0.079383f
C1411 VDD.t104 VSS 0.045109f
C1412 VDD.t10 VSS 0.065453f
C1413 VDD.t113 VSS 0.077172f
C1414 VDD.t288 VSS 0.061191f
C1415 VDD.n60 VSS 0.20297f
C1416 VDD.n61 VSS 0.028256f
C1417 VDD.n62 VSS 0.030799f
C1418 VDD.n63 VSS 0.031942f
C1419 VDD.n64 VSS 0.034152f
C1420 VDD.n65 VSS 0.036128f
C1421 VDD.n66 VSS 0.034475f
C1422 VDD.n67 VSS 0.034441f
C1423 VDD.n68 VSS 0.030226f
C1424 VDD.n69 VSS 0.028068f
C1425 VDD.n70 VSS 0.034252f
C1426 VDD.n71 VSS 0.031942f
C1427 VDD.n72 VSS 0.022319f
C1428 VDD.n73 VSS 0.027693f
C1429 VDD.n74 VSS 0.031942f
C1430 VDD.n75 VSS 0.029317f
C1431 VDD.n76 VSS 0.020695f
C1432 VDD.n77 VSS 0.031942f
C1433 VDD.n78 VSS 0.034252f
C1434 VDD.n79 VSS 0.018134f
C1435 VDD.n80 VSS 0.030369f
C1436 VDD.n81 VSS 0.104621f
C1437 VDD.t29 VSS 0.063905f
C1438 VDD.t6 VSS 0.060367f
C1439 VDD.t296 VSS 0.083806f
C1440 VDD.t318 VSS 0.07872f
C1441 VDD.t126 VSS 0.085133f
C1442 VDD.t93 VSS 0.05904f
C1443 VDD.t98 VSS 0.07872f
C1444 VDD.t286 VSS 0.099063f
C1445 VDD.t181 VSS 0.045109f
C1446 VDD.t2 VSS 0.099063f
C1447 VDD.t25 VSS 0.099285f
C1448 VDD.t139 VSS 0.076449f
C1449 VDD.n82 VSS 0.022845f
C1450 VDD.n83 VSS 0.215558f
C1451 VDD.n84 VSS 0.026348f
C1452 VDD.t187 VSS 0.076363f
C1453 VDD.t78 VSS 0.160382f
C1454 VDD.t100 VSS 0.053902f
C1455 VDD.t74 VSS 0.072901f
C1456 VDD.t70 VSS 0.045508f
C1457 VDD.t27 VSS 0.033282f
C1458 VDD.t116 VSS 0.049484f
C1459 VDD.t199 VSS 0.092341f
C1460 VDD.t183 VSS 0.057437f
C1461 VDD.t153 VSS 0.045066f
C1462 VDD.t251 VSS 0.049484f
C1463 VDD.t155 VSS 0.057437f
C1464 VDD.t151 VSS 0.087481f
C1465 VDD.t204 VSS 0.049484f
C1466 VDD.t149 VSS 0.03159f
C1467 VDD.n94 VSS 0.110506f
C1468 VDD.t171 VSS 0.016347f
C1469 VDD.t138 VSS 0.033579f
C1470 VDD.t51 VSS 0.053019f
C1471 VDD.t233 VSS 0.047717f
C1472 VDD.t130 VSS 0.045066f
C1473 VDD.t173 VSS 0.066052f
C1474 VDD.t298 VSS 0.053902f
C1475 VDD.t235 VSS 0.058541f
C1476 VDD.t68 VSS 0.057437f
C1477 VDD.t203 VSS 0.03888f
C1478 VDD.t53 VSS 0.049484f
C1479 VDD.t72 VSS 0.054786f
C1480 VDD.t169 VSS 0.045066f
C1481 VDD.t76 VSS 0.059204f
C1482 VDD.t66 VSS 0.071575f
C1483 VDD.t55 VSS 0.045066f
C1484 VDD.t80 VSS 0.080854f
C1485 VDD.n95 VSS 0.05946f
C1486 VDD.n97 VSS 0.07635f
C1487 VDD.n98 VSS 0.013402f
C1488 VDD.n99 VSS 0.042269f
C1489 VDD.n100 VSS 0.031334f
C1490 VDD.n101 VSS 0.033863f
C1491 VDD.n102 VSS 0.023862f
C1492 VDD.n103 VSS 0.031631f
C1493 VDD.n104 VSS 0.058048f
C1494 VDD.n105 VSS 0.037311f
C1495 VDD.n106 VSS 0.033112f
C1496 VDD.n107 VSS 0.038664f
C1497 VDD.n108 VSS 0.037258f
C1498 VDD.n109 VSS 0.033155f
C1499 VDD.n110 VSS 0.026353f
C1500 VDD.n111 VSS 0.034072f
C1501 VDD.n112 VSS 0.024692f
C1502 VDD.n113 VSS 0.026687f
C1503 VDD.n114 VSS 0.019167f
C1504 VDD.n117 VSS 0.215659f
C1505 VDD.n118 VSS 0.120425f
C1506 VDD.n119 VSS 0.026348f
C1507 VDD.t49 VSS 0.076363f
C1508 VDD.t267 VSS 0.103387f
C1509 VDD.t224 VSS 0.137407f
C1510 VDD.t82 VSS 0.1405f
C1511 VDD.t19 VSS 0.127024f
C1512 VDD.t246 VSS 0.068927f
C1513 VDD.n126 VSS 0.084555f
C1514 VDD.t86 VSS 0.049042f
C1515 VDD.t0 VSS 0.080412f
C1516 VDD.t4 VSS 0.113769f
C1517 VDD.t88 VSS 0.129012f
C1518 VDD.t18 VSS 0.097422f
C1519 VDD.t31 VSS 0.089248f
C1520 VDD.t132 VSS 0.131663f
C1521 VDD.t33 VSS 0.155963f
C1522 VDD.n127 VSS 0.086411f
C1523 VDD.t134 VSS 0.259792f
C1524 VDD.n128 VSS 0.080667f
C1525 VDD.n129 VSS 0.083864f
C1526 VDD.n130 VSS 0.02608f
C1527 VDD.n131 VSS 0.043514f
C1528 VDD.n132 VSS 0.062247f
C1529 VDD.n133 VSS 0.090658f
C1530 VDD.n134 VSS 0.126497f
C1531 VDD.n135 VSS 0.089224f
C1532 VDD.n136 VSS 0.054943f
C1533 VDD.n137 VSS 0.04188f
C1534 VDD.n138 VSS 0.019167f
C1535 VDD.n139 VSS 0.013085f
C1536 VDD.n141 VSS 0.215659f
C1537 VDD.n142 VSS 0.032616f
C1538 VDD.n143 VSS 0.529173f
C1539 VDD.n144 VSS 0.026348f
C1540 VDD.n145 VSS 0.171639f
C1541 VDD.t261 VSS 0.066815f
C1542 VDD.t47 VSS 0.098968f
C1543 VDD.t16 VSS 0.099189f
C1544 VDD.t290 VSS 0.058983f
C1545 VDD.t244 VSS 0.085051f
C1546 VDD.t21 VSS 0.078644f
C1547 VDD.t60 VSS 0.083725f
C1548 VDD.t111 VSS 0.060309f
C1549 VDD.t96 VSS 0.078644f
C1550 VDD.t272 VSS 0.098968f
C1551 VDD.t45 VSS 0.045066f
C1552 VDD.t12 VSS 0.073343f
C1553 VDD.n146 VSS 0.095026f
C1554 VDD.t84 VSS 0.064064f
C1555 VDD.t58 VSS 0.073343f
C1556 VDD.n147 VSS 0.104526f
C1557 VDD.t114 VSS 0.070913f
C1558 VDD.t62 VSS 0.051914f
C1559 VDD.t274 VSS 0.090132f
C1560 VDD.t89 VSS 0.053019f
C1561 VDD.t64 VSS 0.045066f
C1562 VDD.t294 VSS 0.045066f
C1563 VDD.t276 VSS 0.053019f
C1564 VDD.t8 VSS 0.0581f
C1565 VDD.n150 VSS 0.068471f
C1566 VDD.t278 VSS 0.053163f
C1567 VDD.n151 VSS 0.069951f
C1568 VDD.n152 VSS 0.219068f
C1569 VDD.n153 VSS 0.036104f
C1570 VDD.n154 VSS 0.015075f
C1571 VDD.n155 VSS 0.028404f
C1572 VDD.n156 VSS 0.031567f
C1573 VDD.n157 VSS 0.029348f
C1574 VDD.n158 VSS 0.030334f
C1575 VDD.n159 VSS 0.020121f
C1576 VDD.n160 VSS 0.042269f
C1577 VDD.n161 VSS 0.034379f
C1578 VDD.n162 VSS 0.028322f
C1579 VDD.n163 VSS 0.018095f
C1580 VDD.n164 VSS 0.034157f
C1581 VDD.n165 VSS 0.031855f
C1582 VDD.n166 VSS 0.022639f
C1583 VDD.n167 VSS 0.027246f
C1584 VDD.n168 VSS 0.031855f
C1585 VDD.n169 VSS 0.029612f
C1586 VDD.n170 VSS 0.020272f
C1587 VDD.n171 VSS 0.031855f
C1588 VDD.n172 VSS 0.034157f
C1589 VDD.n173 VSS 0.027995f
C1590 VDD.n174 VSS 0.02116f
C1591 VDD.n175 VSS 0.013085f
C1592 VDD.n177 VSS 0.01137f
C1593 VDD.n179 VSS 0.026392f
C1594 VDD.n181 VSS 0.5353f
C1595 VDD.n182 VSS 0.337617f
C1596 VDD.n183 VSS 5.65783f
C1597 VDD.n184 VSS 0.027798f
C1598 VDD.t280 VSS 0.073714f
C1599 VDD.t36 VSS 0.032909f
C1600 VDD.n185 VSS 0.0719f
C1601 VDD.t253 VSS 0.059477f
C1602 VDD.t42 VSS 0.04524f
C1603 VDD.t300 VSS 0.04524f
C1604 VDD.t136 VSS 0.04524f
C1605 VDD.t258 VSS 0.04524f
C1606 VDD.t257 VSS 0.04524f
C1607 VDD.t259 VSS 0.04524f
C1608 VDD.t260 VSS 0.04524f
C1609 VDD.t44 VSS 0.04524f
C1610 VDD.t14 VSS 0.04524f
C1611 VDD.t106 VSS 0.04524f
C1612 VDD.t15 VSS 0.04524f
C1613 VDD.t284 VSS 0.04524f
C1614 VDD.t37 VSS 0.04524f
C1615 VDD.t308 VSS 0.04524f
C1616 VDD.t102 VSS 0.060083f
C1617 VDD.n186 VSS 0.070546f
C1618 VDD.t103 VSS 0.015288f
C1619 VDD.n188 VSS 0.021218f
C1620 VDD.n189 VSS 0.648587f
C1621 VDD.n190 VSS 0.072942f
C1622 VDD.n191 VSS 0.024032f
C1623 VDD.n192 VSS 0.214671f
C1624 VDD.n193 VSS 0.024032f
C1625 VDD.n194 VSS 0.157507f
C1626 VDD.t254 VSS 0.032909f
C1627 VDD.n195 VSS 0.04969f
C1628 VDD.t283 VSS 0.032909f
C1629 VDD.n196 VSS 0.0719f
C1630 VDD.n197 VSS 0.033006f
C1631 VDD.n198 VSS 0.072779f
C1632 VDD.t282 VSS 0.059477f
C1633 VDD.t137 VSS 0.04524f
C1634 VDD.t285 VSS 0.04524f
C1635 VDD.t35 VSS 0.059477f
C1636 VDD.n199 VSS 0.072779f
C1637 VDD.n200 VSS 0.033006f
C1638 VDD.t281 VSS 0.011082f
C1639 VDD.n201 VSS 0.050108f
C1640 VDD.t307 VSS 0.038748f
C1641 VDD.n202 VSS 0.074374f
C1642 VDD.n203 VSS 0.028818f
C1643 VDD.n204 VSS 0.068663f
C1644 VDD.t303 VSS 0.038748f
C1645 VDD.n205 VSS 0.055484f
C1646 VDD.n206 VSS 0.046977f
C1647 VDD.n207 VSS 0.075839f
C1648 VDD.t302 VSS 0.068658f
C1649 VDD.t304 VSS 0.057481f
C1650 VDD.t107 VSS 0.057481f
C1651 VDD.t306 VSS 0.069245f
C1652 VDD.n208 VSS 0.068748f
C1653 VDD.n209 VSS 0.172389f
C1654 VDD.t123 VSS 0.065403f
C1655 VDD.t122 VSS 0.061008f
C1656 VDD.n215 VSS 0.041107f
C1657 VDD.t121 VSS 0.012419f
C1658 VDD.t311 VSS 0.012419f
C1659 VDD.n217 VSS 0.043721f
C1660 VDD.n218 VSS 0.02442f
C1661 VDD.n223 VSS 0.041107f
C1662 VDD.t119 VSS 0.012419f
C1663 VDD.t186 VSS 0.012419f
C1664 VDD.n225 VSS 0.043721f
C1665 VDD.n226 VSS 0.02442f
C1666 VDD.n231 VSS 0.041107f
C1667 VDD.t125 VSS 0.012419f
C1668 VDD.t191 VSS 0.012419f
C1669 VDD.n233 VSS 0.043721f
C1670 VDD.n234 VSS 0.02442f
C1671 VDD.t129 VSS 0.065833f
C1672 VDD.n240 VSS 0.010214f
C1673 VDD.n242 VSS 0.042777f
C1674 VDD.n243 VSS 0.145691f
C1675 VDD.t128 VSS 0.052139f
C1676 VDD.n244 VSS 0.041107f
C1677 VDD.t124 VSS 0.037308f
C1678 VDD.n245 VSS 0.070815f
C1679 VDD.n257 VSS 0.070815f
C1680 VDD.t190 VSS 0.037308f
C1681 VDD.n258 VSS 0.041107f
C1682 VDD.t118 VSS 0.037308f
C1683 VDD.n259 VSS 0.070815f
C1684 VDD.n271 VSS 0.070815f
C1685 VDD.t185 VSS 0.037308f
C1686 VDD.n272 VSS 0.041107f
C1687 VDD.t120 VSS 0.037308f
C1688 VDD.n273 VSS 0.070815f
C1689 VDD.n286 VSS 0.070815f
C1690 VDD.t310 VSS 0.037308f
C1691 VDD.n287 VSS 0.041107f
C1692 VDD.n288 VSS 0.070815f
C1693 VDD.n291 VSS 0.10548f
C1694 VDD.n292 VSS 0.10519f
C1695 VDD.n294 VSS 0.01751f
C1696 VDD.t144 VSS 0.065902f
C1697 VDD.n310 VSS 0.042845f
C1698 VDD.n311 VSS 0.145927f
C1699 VDD.t143 VSS 0.05226f
C1700 VDD.n314 VSS 0.070946f
C1701 VDD.t147 VSS 0.037376f
C1702 VDD.n318 VSS 0.070946f
C1703 VDD.t145 VSS 0.037376f
C1704 VDD.n322 VSS 0.070946f
C1705 VDD.t206 VSS 0.037376f
C1706 VDD.t211 VSS 0.065472f
C1707 VDD.n326 VSS 0.10527f
C1708 VDD.n329 VSS 0.105656f
C1709 VDD.t210 VSS 0.061151f
C1710 VDD.n330 VSS 0.070946f
C1711 VDD.n331 VSS 0.041183f
C1712 VDD.t110 VSS 0.012419f
C1713 VDD.t207 VSS 0.012419f
C1714 VDD.n333 VSS 0.043777f
C1715 VDD.n334 VSS 0.024421f
C1716 VDD.n339 VSS 0.041183f
C1717 VDD.t109 VSS 0.037376f
C1718 VDD.n340 VSS 0.070946f
C1719 VDD.n341 VSS 0.041183f
C1720 VDD.t198 VSS 0.012419f
C1721 VDD.t146 VSS 0.012419f
C1722 VDD.n343 VSS 0.043777f
C1723 VDD.n344 VSS 0.024421f
C1724 VDD.n349 VSS 0.041183f
C1725 VDD.t197 VSS 0.037376f
C1726 VDD.n350 VSS 0.070946f
C1727 VDD.n351 VSS 0.041183f
C1728 VDD.t209 VSS 0.012419f
C1729 VDD.t148 VSS 0.012419f
C1730 VDD.n353 VSS 0.043777f
C1731 VDD.n354 VSS 0.024421f
C1732 VDD.n359 VSS 0.041183f
C1733 VDD.t208 VSS 0.037376f
C1734 VDD.n360 VSS 0.070946f
C1735 VDD.n361 VSS 0.041183f
C1736 VDD.n365 VSS 0.666268f
C1737 VDD.n366 VSS 5.27642f
C1738 VDD.n367 VSS 1.84975f
C1739 VDD.n368 VSS 2.63548f
C1740 VDD.n369 VSS 0.937979f
C1741 VDD.t229 VSS 0.0853f
C1742 VDD.n372 VSS 0.056987f
C1743 VDD.t215 VSS 0.118367f
C1744 VDD.n373 VSS 0.118192f
C1745 VDD.n374 VSS 0.010102f
C1746 VDD.n375 VSS 0.084411f
C1747 VDD.n376 VSS 0.38652f
C1748 VDD.t220 VSS 0.0853f
C1749 VDD.n379 VSS 0.056987f
C1750 VDD.t28 VSS 0.118367f
C1751 VDD.n380 VSS 0.118192f
C1752 VDD.n381 VSS 0.010102f
C1753 VDD.n382 VSS 0.084411f
C1754 VDD.n383 VSS 0.46741f
C1755 VDD.t237 VSS 0.0853f
C1756 VDD.n386 VSS 0.056987f
C1757 VDD.t249 VSS 0.118367f
C1758 VDD.n387 VSS 0.118192f
C1759 VDD.n388 VSS 0.010102f
C1760 VDD.n389 VSS 0.084411f
C1761 VDD.n390 VSS 0.46741f
C1762 VDD.t222 VSS 0.0853f
C1763 VDD.n393 VSS 0.056987f
C1764 VDD.t41 VSS 0.118367f
C1765 VDD.n394 VSS 0.118192f
C1766 VDD.n395 VSS 0.010102f
C1767 VDD.n396 VSS 0.084411f
C1768 VDD.n397 VSS 0.46741f
C1769 VDD.t227 VSS 0.0853f
C1770 VDD.n400 VSS 0.056987f
C1771 VDD.t95 VSS 0.118367f
C1772 VDD.n401 VSS 0.118192f
C1773 VDD.n402 VSS 0.010102f
C1774 VDD.n403 VSS 0.084411f
C1775 VDD.n404 VSS 0.46741f
C1776 VDD.t231 VSS 0.0853f
C1777 VDD.n407 VSS 0.056987f
C1778 VDD.t189 VSS 0.118367f
C1779 VDD.n408 VSS 0.118192f
C1780 VDD.n409 VSS 0.010102f
C1781 VDD.n410 VSS 0.084411f
C1782 VDD.n411 VSS 0.46741f
C1783 VDD.n412 VSS 0.73398f
C1784 VDD.t218 VSS 0.0853f
C1785 VDD.n413 VSS 0.090631f
C1786 VDD.t265 VSS 0.0853f
C1787 VDD.n414 VSS 0.095369f
C1788 VDD.n415 VSS 0.056123f
C1789 VDD.n416 VSS 0.626949f
C1790 VDD.n417 VSS 5.28484f
.ends

