* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP DEBUG VDD PLL_FREERUN VSS PLL_CLK_OUT PLL_DISABLE PLL_REF_CLK PLL_VCTRL
X0 a_23444_3994 a_22864_4398 VSS.t327 VSS.t326 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 VDD.t182 a_22948_2038 a_22864_2486 VDD.t181 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X2 a_23099_4907 a_23011_4951 VSS.t252 VSS.t251 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_24355_n1338.t27 a_23423_n1258 VSS.t250 VSS.t249 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4 a_24355_n1338.t36 a_27899_438.t13 PLL_CLK_OUT.t28 VSS.t254 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X5 a_5840_15093.t9 a_5840_7613.t0 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X6 VSS.t85 a_23455_217 a_23407_261 VSS.t40 nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X7 a_22864_4398 a_22948_3950 a_22884_3994 VSS.t153 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X8 a_24355_n1338.t37 a_27899_438.t14 PLL_CLK_OUT.t27 VSS.t255 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X9 PLL_CLK_OUT.t26 a_27899_438.t15 a_24355_n1338.t38 VSS.t256 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X10 VDD.t329 a_22388_2038.t2 a_22304_2486 VDD.t328 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X11 DEBUG.t25 PLL_FREERUN.t0 PLL_VCTRL.t15 VSS.t259 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X12 a_n2908_12013 a_1220_12453 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X13 VSS.t61 a_31031_1644 a_30943_1688 VSS.t60 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X14 a_24891_4907 a_24803_4951 VSS.t348 VSS.t347 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X15 PLL_CLK_OUT.t34 PLL_DISABLE.t0 a_24355_n1338.t47 VDD.t327 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X16 a_5840_15093.t9 a_5840_7613.t0 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X17 a_n15085_2072.t19 PLL_FREERUN.t1 DEBUG.t29 VDD.t266 pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.33u
X18 a_22539_3430 a_22451_3522 VDD.t176 VDD.t175 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X19 a_n558_2704.t1 a_11009_2840 a_14657_n1138 VSS.t196 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X20 DEBUG.t24 PLL_FREERUN.t2 PLL_VCTRL.t14 VSS.t268 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X21 a_n15085_2072.t32 a_n17351_68.t2 DEBUG.t62 VSS.t267 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X22 a_22203_n358.t3 a_21855_n1258 VSS.t57 VSS.t56 nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
X23 VSS.t124 a_23455_1567 a_23407_1611 VSS.t123 nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X24 a_n15085_2072.t41 VSS.t188 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X25 a_21855_4398 a_21755_4018 VSS.t178 VSS.t177 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X26 PLL_VCTRL.t31 a_n17351_68.t3 DEBUG.t63 VDD.t264 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X27 PLL_VCTRL.t32 a_n17351_68.t4 DEBUG.t64 VDD.t265 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X28 DEBUG.t52 a_n17351_68.t5 PLL_VCTRL.t24 VDD.t183 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X29 a_25265_7733 a_24755_6933 a_5840_15093.t3 VDD.t128 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X30 VSS.t248 a_23423_n1258 a_24355_n1338.t26 VSS.t247 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X31 a_22203_n358.t2 a_21855_n1258 VSS.t55 VSS.t54 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X32 DEBUG.t53 a_n17351_68.t6 PLL_VCTRL.t25 VDD.t184 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X33 VSS.t211 a_n4208_n141.t3 a_n671_n1138 VSS.t210 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X34 VDD.t201 a_n8471_219.t5 a_3149_2840 VDD.t200 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X35 a_21755_1082 a_24383_1567 VSS.t342 VSS.t341 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X36 PLL_VCTRL.t26 a_n17351_68.t7 DEBUG.t54 VDD.t185 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X37 a_27491_1710 PLL_REF_CLK.t0 VSS.t147 VSS.t146 nfet_06v0 ad=0.1584p pd=1.6u as=0.151p ps=1.185u w=0.36u l=0.6u
X38 a_24355_n1338.t8 PLL_DISABLE.t1 PLL_CLK_OUT.t3 VDD.t112 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X39 VDD.t83 a_23620_8319.t3 a_23691_7733 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.52p ps=2.52u w=2u l=0.33u
X40 DEBUG.t28 PLL_FREERUN.t3 a_n15085_2072.t18 VDD.t267 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X41 VSS.t41 a_23455_n345 a_23407_n301 VSS.t40 nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X42 VSS.t143 a_n8537_n1530.t4 a_n8659_n1230 VSS.t142 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X43 a_22987_3430 a_22899_3522 VDD.t241 VDD.t240 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X44 a_25675_477 a_25587_574 VSS.t30 VSS.t29 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X45 VDD.t209 a_22203_n358.t8 a_22115_253.t1 VDD.t208 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X46 a_7177_2840 a_3345_2840 a_6981_2840 VDD.t80 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X47 VDD.t77 a_23508_2038 a_22948_2038 VDD.t76 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X48 a_27014_14933 a_24866_11400 VSS.t68 ppolyf_u r_width=0.8u r_length=22u
X49 a_n15085_2072.t42 VSS.t189 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X50 DEBUG.t68 a_n17351_68.t8 PLL_VCTRL.t33 VDD.t272 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X51 VDD.t47 a_21855_n1258 a_22203_n358.t7 VDD.t46 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X52 a_22948_3950 a_23508_2038 a_23444_3994 VSS.t84 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X53 a_5840_15093.t9 a_5840_7613.t0 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X54 a_26795_6933 a_n8537_93.t3 a_25265_6933 VSS.t98 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X55 PLL_VCTRL.t34 a_n17351_68.t9 DEBUG.t69 VDD.t273 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X56 a_24355_n1338.t41 a_27899_438.t16 PLL_CLK_OUT.t25 VSS.t285 nfet_03v3 ad=0.65p pd=3.3u as=0.26p ps=1.52u w=1u l=0.33u
X57 a_1220_13333 a_5840_13333 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X58 PLL_CLK_OUT.t24 a_27899_438.t17 a_24355_n1338.t42 VSS.t286 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X59 PLL_CLK_OUT.t4 PLL_DISABLE.t2 a_24355_n1338.t9 VDD.t113 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X60 a_24355_n1338.t43 a_27899_438.t18 PLL_CLK_OUT.t23 VSS.t287 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X61 a_n15085_2072.t36 a_n17351_68.t10 DEBUG.t70 VSS.t284 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X62 VDD.t257 a_21394_11355.t16 a_21394_11355.t17 VDD.t256 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X63 a_24383_217 a_24090_629 VDD.t116 VDD.t115 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X64 DEBUG.t77 a_n17351_68.t11 PLL_VCTRL.t38 VDD.t342 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X65 a_1712_14653 a_5840_15093.t4 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X66 VSS.t313 a_16431_6193 VSS.t183 ppolyf_u r_width=0.8u r_length=0.13m
X67 a_26049_6873 a_25369_6873 VDD.t277 VDD.t276 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X68 a_23407_1611 a_22527_1197 a_23083_1611 VSS.t67 nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X69 a_21643_3430 a_21555_3522 VDD.t52 VDD.t51 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X70 a_n8471_219.t0 a_n8537_93.t4 a_n8659_n1230 VSS.t99 nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.33u
X71 PLL_CLK_OUT.t5 PLL_DISABLE.t3 a_24355_n1338.t10 VDD.t114 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X72 a_22864_4398 a_22304_4398 VDD.t28 VDD.t27 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X73 a_21506_13215.t9 a_21394_11355.t18 VDD.t259 VDD.t258 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X74 a_23083_1611 a_22963_1518 a_22915_1611 VSS.t308 nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X75 DEBUG.t27 PLL_FREERUN.t4 a_n15085_2072.t17 VDD.t194 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X76 a_n2908_11133 a_1220_11573 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X77 VSS.t346 a_24675_7463 a_24755_6933 VSS.t345 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X78 a_22304_4398 a_21855_4398 VDD.t317 VDD.t316 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X79 PLL_VCTRL.t39 a_n17351_68.t12 DEBUG.t78 VDD.t343 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X80 DEBUG.t79 a_n17351_68.t13 a_n15085_2072.t40 VSS.t335 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X81 a_24355_n1338.t35 a_23423_n1258 VDD.t236 VDD.t235 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X82 VDD.t203 a_n8471_219.t6 a_18477_2840 VDD.t202 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X83 VDD.t220 a_22864_2486 a_22388_2038.t1 VDD.t219 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X84 VDD.t234 a_23423_n1258 a_24355_n1338.t34 VDD.t233 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X85 DEBUG.t74 a_n17351_68.t14 PLL_VCTRL.t35 VDD.t324 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X86 VSS.t246 a_23423_n1258 a_24355_n1338.t25 VSS.t245 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X87 a_22959_n669 a_22527_n715 VDD.t50 VDD.t49 pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X88 VSS.t111 a_25675_n394 a_25587_n302 VSS.t29 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X89 a_23083_261 a_22963_217 a_22915_261 VSS.t14 nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X90 VDD.t247 a_21394_11355.t19 a_21506_13215.t8 VDD.t246 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X91 a_23407_n301 a_22527_n715 a_23083_n301 VSS.t59 nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X92 a_21855_1126 a_21755_1082 VSS.t301 VSS.t299 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X93 a_21855_n1258 a_n558_2704.t2 VSS.t312 VSS.t311 nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X94 PLL_VCTRL.t36 a_n17351_68.t15 DEBUG.t75 VDD.t325 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X95 VSS.t145 a_n8537_n1530.t5 a_21891_6933 VSS.t144 nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.33u
X96 a_22959_1243 a_22527_1197 VDD.t58 VDD.t57 pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X97 a_n15085_2072.t43 VSS.t191 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X98 PLL_VCTRL.t37 a_n17351_68.t16 DEBUG.t76 VDD.t326 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X99 a_25265_7733 a_22941_7733.t3 a_25095_7733 VDD.t64 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X100 a_24355_n1338.t46 PLL_DISABLE.t4 PLL_CLK_OUT.t33 VDD.t283 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X101 a_5840_15093.t9 a_5840_7613.t0 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X102 a_23083_n301 a_21855_1126 a_22915_n301 VSS.t14 nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X103 DEBUG.t55 a_n17351_68.t17 PLL_VCTRL.t27 VDD.t196 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X104 VSS.t193 a_n8537_n1530.t6 a_n8659_n1230 VSS.t192 nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.33u
X105 a_n15085_2072.t29 a_n17351_68.t18 DEBUG.t56 VSS.t224 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X106 a_22941_7733.t2 a_n8537_93.t5 a_22955_6933 VSS.t138 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X107 a_n15085_2072.t16 PLL_FREERUN.t5 DEBUG.t26 VDD.t195 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X108 a_24383_n345 a_24090_n669 VDD.t30 VDD.t29 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X109 a_23427_629 a_22115_253.t2 a_23083_261 VDD.t102 pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X110 a_21755_1082 a_24383_1567 VDD.t347 VDD.t92 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X111 a_22527_1197 a_22115_1610.t2 VSS.t20 VSS.t19 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X112 VDD.t210 a_22203_n358.t9 a_22115_1610.t1 VDD.t208 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X113 a_21855_n1258 a_n558_2704.t3 VDD.t172 VDD.t171 pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X114 PLL_CLK_OUT.t22 a_27899_438.t19 a_24355_n1338.t11 VSS.t165 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X115 a_21506_13215.t7 a_21394_11355.t20 VDD.t249 VDD.t248 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X116 a_24355_n1338.t12 a_27899_438.t20 PLL_CLK_OUT.t21 VSS.t166 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X117 PLL_CLK_OUT.t20 a_27899_438.t21 a_24355_n1338.t13 VSS.t167 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X118 DEBUG.t23 PLL_FREERUN.t6 PLL_VCTRL.t7 VSS.t223 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X119 a_24355_n1338.t24 a_23423_n1258 VSS.t244 VSS.t243 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X120 a_22527_574 a_22115_253.t3 VDD.t104 VDD.t103 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X121 a_23083_n301 a_21855_1126 a_22959_n669 VDD.t10 pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X122 a_26115_6933 a_26049_6873 a_25265_6933 VSS.t115 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X123 VSS.t91 a_22091_3430 a_22003_3522 VSS.t90 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X124 a_23407_261 a_22527_574 a_23083_261 VSS.t59 nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X125 DEBUG.t39 PLL_FREERUN.t7 a_n15085_2072.t15 VDD.t198 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X126 a_23083_1611 a_22963_1518 a_22959_1243 VDD.t59 pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X127 a_22915_1611 a_22115_1610.t3 VSS.t119 VSS.t118 nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X128 a_22948_3950 a_22864_4398 VDD.t335 VDD.t334 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X129 a_22203_n358.t6 a_21855_n1258 VDD.t45 VDD.t44 pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X130 a_23435_3430 a_23347_3522 VDD.t292 VDD.t291 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D0 PLL_DISABLE.t5 VDD.t284 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X131 PLL_VCTRL.t28 a_n17351_68.t19 DEBUG.t57 VDD.t197 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X132 DEBUG.t58 a_n17351_68.t20 a_n15085_2072.t30 VSS.t257 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X133 VDD.t218 a_22864_2486 a_23508_2038 VDD.t217 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X134 a_24207_4398 a_22304_4398 VSS.t35 VSS.t34 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X135 a_23455_217 a_23083_261 VSS.t13 VSS.t12 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X136 VDD.t243 a_n8471_219.t3 a_n8471_219.t4 VDD.t242 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X137 a_25265_7733 a_24675_7463 a_26115_6933 VDD.t355 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X138 a_23423_n1258 a_22203_n358.t10 VSS.t230 VSS.t229 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X139 PLL_VCTRL.t6 PLL_FREERUN.t8 DEBUG.t22 VSS.t225 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X140 a_22203_n358.t5 a_21855_n1258 VDD.t43 VDD.t42 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X141 a_24355_n1338.t33 a_23423_n1258 VDD.t232 VDD.t231 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X142 VDD.t345 a_25675_477 a_25587_574 VDD.t318 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X143 a_23423_n1258 a_22203_n358.t11 VSS.t202 VSS.t201 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X144 a_22915_n301 a_22115_n302.t2 VSS.t298 VSS.t151 nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X145 VDD.t79 a_23455_217 a_23427_629 VDD.t78 pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X146 a_n15085_2072.t44 VSS.t319 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X147 a_23691_7733 a_23620_8319.t4 VDD.t85 VDD.t84 pfet_03v3 ad=0.52p pd=2.52u as=1.3p ps=5.3u w=2u l=0.33u
X148 a_n2908_7613 VSS.t160 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X149 VSS.t195 a_n8537_n1530.t7 a_22955_6933 VSS.t194 nfet_03v3 ad=0.4p pd=1.8u as=0.26p ps=1.52u w=1u l=0.33u
X150 a_n15085_2072.t14 PLL_FREERUN.t9 DEBUG.t38 VDD.t199 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X151 a_22388_3950.t0 a_23508_2038 VDD.t75 VDD.t74 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X152 a_n2908_10253 a_1220_10693 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X153 a_23883_3430 a_23795_3522 VDD.t3 VDD.t2 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X154 a_24655_4398 a_24207_4398 VSS.t24 VSS.t23 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X155 a_n2908_9373 a_1220_8933 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X156 VDD.t314 a_21755_4907 a_21667_4951 VDD.t313 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X157 PLL_CLK_OUT.t19 a_27899_438.t22 a_24355_n1338.t3 VSS.t135 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X158 a_21855_4398 a_21755_4018 VDD.t124 VDD.t123 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X159 a_22388_3950.t0 a_24655_4398 VDD.t66 VDD.t65 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X160 DEBUG.t21 PLL_FREERUN.t10 PLL_VCTRL.t17 VSS.t317 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X161 a_21755_477 a_21667_574 VSS.t76 VSS.t43 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X162 a_11009_2840 a_7177_2840 a_10813_2840 VDD.t69 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X163 VDD.t166 a_n8471_219.t7 a_n683_2840 VDD.t165 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X164 a_24675_7463 a_22388_3950.t2 VSS.t73 VSS.t72 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X165 PLL_VCTRL.t29 a_n17351_68.t21 DEBUG.t59 VDD.t238 pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.33u
X166 a_n15085_2072.t31 a_n17351_68.t22 DEBUG.t60 VSS.t258 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X167 a_26115_6933 a_26049_6873 a_25265_6933 VSS.t114 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X168 VDD.t22 a_27491_1710 a_21755_4018 VDD.t21 pfet_06v0 ad=0.458p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
X169 a_25150_3994 a_24655_4398 VSS.t78 VSS.t77 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X170 a_22304_4398 a_22388_3950.t3 a_22324_3994 VSS.t49 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X171 DEBUG.t37 PLL_FREERUN.t11 a_n15085_2072.t13 VDD.t323 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X172 VSS.t53 a_21855_n1258 a_22203_n358.t1 VSS.t52 nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X173 DEBUG.t20 PLL_FREERUN.t12 PLL_VCTRL.t16 VSS.t318 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X174 a_27899_438.t10 PLL_DISABLE.t6 VDD.t286 VDD.t285 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X175 a_21506_13215.t6 a_21394_11355.t21 VDD.t251 VDD.t250 pfet_03v3 ad=1.456p pd=6.12u as=3.64p ps=12.5u w=5.6u l=0.56u
X176 VSS.t204 a_22203_n358.t12 a_22115_1610.t0 VSS.t203 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X177 a_22963_217 a_24383_n345 VDD.t7 VDD.t6 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X178 a_25265_7733 a_24675_7463 a_26115_6933 VDD.t354 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X179 a_22388_2038.t0 a_23508_2038 a_25334_2082 VSS.t83 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X180 a_23620_8319.t2 a_n8537_93.t6 a_23691_6933 VSS.t139 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X181 VDD.t189 a_21394_11355.t22 a_21506_13215.t5 VDD.t188 pfet_03v3 ad=3.64p pd=12.5u as=1.456p ps=6.12u w=5.6u l=0.56u
X182 a_1712_7613 a_5840_7613.t1 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X183 VDD.t340 a_22941_7733.t0 a_22941_7733.t1 VDD.t339 pfet_03v3 ad=1.072p pd=5.3u as=1.072p ps=5.3u w=0.8u l=0.33u
X184 a_31479_1644 a_31391_1688 VDD.t39 VDD.t38 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X185 VDD.t95 a_24383_217 a_24375_629 VDD.t94 pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X186 a_24355_n1338.t44 PLL_DISABLE.t7 PLL_CLK_OUT.t31 VDD.t279 pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.33u
X187 DEBUG.t49 a_n17351_68.t23 a_n15085_2072.t26 VSS.t168 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X188 VDD.t97 a_n558_2704.t4 a_21855_n1258 VDD.t96 pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X189 a_1712_9373 a_5840_8933 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X190 a_23691_7733 a_22941_7733.t4 a_23620_8319.t1 VDD.t100 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X191 a_21755_4018 a_27491_1710 VSS.t28 VSS.t27 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X192 a_27899_438.t9 PLL_DISABLE.t8 VDD.t281 VDD.t280 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X193 a_24355_n1338.t45 PLL_DISABLE.t9 PLL_CLK_OUT.t32 VDD.t282 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X194 a_21891_6933 a_n8537_n1530.t8 VSS.t101 VSS.t100 nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.33u
X195 a_1712_11133 a_5840_11573 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X196 a_n2908_14213 a_1220_14653 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X197 a_24755_6933 a_24675_7463 VDD.t353 VDD.t352 pfet_03v3 ad=0.52p pd=2.52u as=1.3p ps=5.3u w=2u l=0.33u
X198 a_22915_261 a_22115_253.t4 VSS.t152 VSS.t151 nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X199 a_24090_629 a_22115_253.t5 a_23455_217 VDD.t86 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X200 a_5840_15093.t9 a_5840_7613.t0 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X201 a_27899_438.t5 PLL_DISABLE.t10 VDD.t364 VDD.t363 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X202 a_n15085_2072.t27 a_n17351_68.t24 DEBUG.t50 VSS.t169 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X203 VDD.t191 a_21394_11355.t23 a_21506_13215.t4 VDD.t190 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X204 DEBUG.t5 PLL_FREERUN.t13 a_n15085_2072.t12 VDD.t320 pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.33u
X205 a_n15085_2072.t11 PLL_FREERUN.t14 DEBUG.t4 VDD.t321 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X206 VSS.t110 a_n8537_93.t1 a_n8537_93.t2 VSS.t109 nfet_03v3 ad=0.496p pd=3.22u as=0.496p ps=3.22u w=0.4u l=0.33u
X207 a_24355_n1338.t4 a_27899_438.t23 PLL_CLK_OUT.t18 VSS.t136 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X208 VDD.t310 a_23547_4907 a_23459_4951 VDD.t309 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X209 PLL_CLK_OUT.t17 a_27899_438.t24 a_24355_n1338.t5 VSS.t137 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X210 VSS.t206 a_22203_n358.t13 a_23423_n1258 VSS.t205 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X211 a_27814_14933 a_27414_10401 VSS.t42 ppolyf_u r_width=0.8u r_length=22u
X212 a_25104_3522 a_22304_4398 a_24900_3522 VSS.t33 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X213 a_3345_2840 a_n487_2840 a_3149_2840 VDD.t81 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X214 a_5840_15093.t9 a_5840_7613.t0 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X215 a_25334_3994 a_22864_4398 a_25150_3994 VSS.t325 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X216 a_22884_2082 a_22304_2486 VSS.t307 VSS.t306 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X217 VDD.t294 a_23620_8319.t5 a_26795_7733 VDD.t293 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X218 a_22527_574 a_22115_253.t6 VSS.t107 VSS.t106 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X219 PLL_CLK_OUT.t38 PLL_DISABLE.t11 a_24355_n1338.t54 VDD.t365 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X220 a_n2908_8493 a_1220_8053 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X221 a_25265_6933 a_25369_6873 a_5840_15093.t8 VSS.t295 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X222 a_n15085_2072.t45 VSS.t188 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X223 a_22324_2082 a_21855_2486 VSS.t70 VSS.t69 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X224 a_7177_2840 a_3345_2840 a_6993_n1138 VSS.t92 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X225 a_21755_4018 a_27491_1710 VDD.t20 VDD.t19 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X226 a_n487_2840 a_n558_2704.t5 a_n671_n1138 VSS.t266 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X227 a_5840_15093.t9 a_5840_7613.t0 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X228 a_21394_11355.t15 a_21394_11355.t14 VDD.t157 VDD.t156 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X229 a_23455_n345 a_23083_n301 VDD.t68 VDD.t67 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X230 a_24335_261 a_22115_253.t7 a_24090_629 VSS.t108 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X231 VDD.t357 a_22203_4907 a_22115_4951 VDD.t356 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X232 a_5840_15093.t2 a_24755_6933 a_25265_7733 VDD.t127 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X233 a_22527_n715 a_22115_n302.t3 VDD.t290 VDD.t289 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X234 VDD.t12 a_23995_4907 a_23907_4951 VDD.t11 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X235 a_23455_1567 a_23083_1611 VDD.t31 VDD.t8 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X236 a_n4208_n141.t2 a_n8471_219.t8 VDD.t168 VDD.t167 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X237 a_n15085_2072.t10 PLL_FREERUN.t15 DEBUG.t3 VDD.t322 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X238 a_24355_n1338.t55 PLL_DISABLE.t12 PLL_CLK_OUT.t39 VDD.t366 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X239 a_27899_438.t12 PLL_DISABLE.t13 VDD.t360 VDD.t359 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X240 a_24355_n1338.t32 a_23423_n1258 VDD.t230 VDD.t229 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X241 VSS.t242 a_23423_n1258 a_24355_n1338.t23 VSS.t241 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X242 a_23455_217 a_23083_261 VDD.t9 VDD.t8 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X243 VDD.t1 a_21755_477 a_21667_574 VDD.t0 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X244 a_22955_6933 a_n8537_n1530.t9 VSS.t103 VSS.t102 nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.33u
X245 a_n15085_2072.t46 VSS.t189 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X246 a_1712_8493 a_5840_8053 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X247 a_24355_n1338.t17 a_27899_438.t25 PLL_CLK_OUT.t16 VSS.t219 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X248 a_24207_4398 a_22304_4398 VDD.t26 VDD.t25 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X249 VSS.t16 a_25675_1518 a_25587_1610 VSS.t15 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X250 a_21855_2486 a_21755_1082 VSS.t300 VSS.t299 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X251 VDD.t130 a_22651_4907 a_22563_4951 VDD.t129 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X252 a_23444_2082 a_22864_2486 VSS.t234 VSS.t233 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X253 VDD.t302 a_25339_4907 a_25251_4951 VDD.t301 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X254 a_18673_2840 a_n558_2704.t6 a_18477_2840 VDD.t162 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X255 a_1712_10253 a_5840_10693 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X256 a_24383_217 a_24090_629 VSS.t161 VSS.t36 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X257 a_n2908_13333 a_1220_13773 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X258 a_25265_6933 a_25369_6873 a_5840_15093.t7 VSS.t294 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X259 DEBUG.t51 a_n17351_68.t25 a_n15085_2072.t28 VSS.t170 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X260 VDD.t41 a_21855_n1258 a_22203_n358.t4 VDD.t40 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X261 VDD.t33 a_23455_n345 a_23427_n669 VDD.t32 pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X262 PLL_VCTRL.t1 PLL_FREERUN.t16 DEBUG.t19 VSS.t148 nfet_03v3 ad=0.26p pd=1.52u as=0.65p ps=3.3u w=1u l=0.33u
X263 a_21855_1126 a_21755_1082 VDD.t300 VDD.t299 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X264 a_22864_2486 a_22948_2038 a_22884_2082 VSS.t216 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X265 VSS.t87 a_n8537_n1530.t10 a_23691_6933 VSS.t86 nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.33u
X266 PLL_CLK_OUT.t36 PLL_DISABLE.t14 a_24355_n1338.t52 VDD.t361 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X267 VDD.t91 a_23455_1567 a_23427_1243 VDD.t78 pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X268 a_23508_2038 a_22304_2486 VDD.t308 VDD.t307 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X269 a_n8471_219.t2 DEBUG.t80 a_n9701_6193 VSS.t198 nfet_03v3 ad=0.488p pd=2.82u as=0.488p ps=2.82u w=0.8u l=0.33u
X270 PLL_VCTRL.t0 PLL_FREERUN.t17 DEBUG.t18 VSS.t149 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X271 a_18673_2840 a_n558_2704.t7 a_18489_n1138 VSS.t226 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X272 a_24655_4398 a_24207_4398 VDD.t16 VDD.t15 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X273 VDD.t159 a_22203_n358.t14 a_23423_n1258 VDD.t158 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
D1 VSS.t63 VSS.t62 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X274 a_n15085_2072.t9 PLL_FREERUN.t18 DEBUG.t2 VDD.t106 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X275 a_n2908_12013 a_1220_11573 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X276 a_24383_1567 a_24090_1243 VSS.t172 VSS.t171 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X277 a_24675_7463 a_22388_3950.t4 VDD.t37 VDD.t36 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X278 PLL_VCTRL.t13 PLL_FREERUN.t19 DEBUG.t17 VSS.t273 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X279 a_23508_2038 a_22864_4398 a_25104_3522 VSS.t324 nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X280 a_25095_7733 a_23620_8319.t6 VDD.t296 VDD.t295 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X281 a_23455_1567 a_23083_1611 VSS.t39 VSS.t38 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X282 a_22091_3430 a_22003_3522 VDD.t18 VDD.t17 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X283 a_24866_11400 a_21506_13215.t10 a_21394_11355.t0 VSS.t2 nfet_03v3 ad=3.416p pd=12.42u as=1.456p ps=6.12u w=5.6u l=0.56u
X284 DEBUG.t16 PLL_FREERUN.t20 PLL_VCTRL.t12 VSS.t274 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X285 a_26049_6873 a_25369_6873 VSS.t293 VSS.t292 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X286 a_22959_629 a_22527_574 VDD.t90 VDD.t57 pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X287 a_22864_2486 a_22304_2486 VDD.t306 VDD.t305 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X288 VSS.t213 a_n4208_n141.t4 a_18489_n1138 VSS.t212 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X289 a_31031_1644 a_30943_1688 VDD.t263 VDD.t262 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X290 a_24383_n345 a_24090_n669 VSS.t37 VSS.t36 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X291 DEBUG.t65 a_n17351_68.t26 a_n15085_2072.t33 VSS.t270 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X292 VDD.t228 a_23423_n1258 a_24355_n1338.t31 VDD.t227 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X293 a_27491_1710 PLL_REF_CLK.t1 VDD.t146 VDD.t145 pfet_06v0 ad=0.4488p pd=2.92u as=0.458p ps=2.02u w=1.02u l=0.5u
X294 a_22304_2486 a_21855_2486 VDD.t61 VDD.t60 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X295 VDD.t35 a_24443_4907 a_24355_4951 VDD.t34 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X296 DEBUG.t15 PLL_FREERUN.t21 PLL_VCTRL.t3 VSS.t275 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X297 a_1712_14653 a_5840_14213 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X298 VDD.t275 a_25369_6873 a_26049_6873 VDD.t274 pfet_03v3 ad=1.3p pd=5.3u as=0.52p ps=2.52u w=2u l=0.33u
X299 a_22948_2038 a_23508_2038 a_23444_2082 VSS.t82 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X300 VDD.t333 a_22864_4398 a_23508_2038 VDD.t332 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X301 a_5840_15093.t9 a_5840_7613.t0 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X302 a_23455_n345 a_23083_n301 VSS.t79 VSS.t12 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X303 a_24383_1567 a_24090_1243 VDD.t119 VDD.t115 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X304 DEBUG.t14 PLL_FREERUN.t22 PLL_VCTRL.t2 VSS.t150 nfet_03v3 ad=0.65p pd=3.3u as=0.26p ps=1.52u w=1u l=0.33u
X305 a_25265_6933 a_n8537_93.t7 a_25095_6933 VSS.t140 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X306 a_n15085_2072.t8 PLL_FREERUN.t23 DEBUG.t1 VDD.t107 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X307 a_n2908_9373 a_1220_9813 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X308 a_24355_n1338.t53 PLL_DISABLE.t15 PLL_CLK_OUT.t37 VDD.t362 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X309 VDD.t261 a_23099_4907 a_23011_4951 VDD.t260 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X310 VDD.t121 a_21755_n830 a_21667_n786 VDD.t120 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X311 a_n487_2840 a_n558_2704.t8 a_n683_2840 VDD.t131 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X312 a_5840_15093.t1 a_24755_6933 a_25265_7733 VDD.t126 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X313 a_24355_n1338.t39 PLL_DISABLE.t16 PLL_CLK_OUT.t29 VDD.t268 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X314 VDD.t312 a_24891_4907 a_24803_4951 VDD.t311 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X315 a_21394_11355.t13 a_21394_11355.t12 VDD.t214 VDD.t213 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X316 a_n15085_2072.t34 a_n17351_68.t27 DEBUG.t66 VSS.t271 nfet_03v3 ad=0.26p pd=1.52u as=0.65p ps=3.3u w=1u l=0.33u
X317 a_22955_6933 a_n8537_93.t8 a_22941_7733.t2 VSS.t141 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X318 DEBUG.t0 PLL_FREERUN.t24 a_n15085_2072.t7 VDD.t108 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X319 VDD.t5 a_24383_n345 a_24375_n669 VDD.t4 pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X320 VDD.t346 a_24383_1567 a_24375_1243 VDD.t94 pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X321 a_24375_629 a_22527_574 a_24090_629 VDD.t56 pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X322 a_22948_2038 a_22864_2486 VDD.t216 VDD.t215 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X323 a_n2908_11133 a_1220_10693 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X324 PLL_CLK_OUT.t15 a_27899_438.t26 a_24355_n1338.t18 VSS.t220 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X325 a_24207_2486 a_22304_2486 VSS.t305 VSS.t304 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X326 a_n15085_2072.t47 VSS.t190 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X327 VDD.t212 a_21394_11355.t10 a_21394_11355.t11 VDD.t211 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X328 a_25265_6933 a_26049_6873 a_26115_6933 VSS.t113 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X329 PLL_CLK_OUT.t30 PLL_DISABLE.t17 a_24355_n1338.t40 VDD.t269 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X330 a_22963_1518 a_24383_217 VSS.t130 VSS.t10 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X331 a_1712_9373 a_5840_9813 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X332 a_n15085_2072.t6 PLL_FREERUN.t25 DEBUG.t36 VDD.t186 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X333 VDD.t110 a_22948_3950 a_22864_4398 VDD.t109 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X334 VSS.t3 a_24866_11400 a_21506_13215.t1 VSS.t2 nfet_03v3 ad=3.416p pd=12.42u as=1.456p ps=6.12u w=5.6u l=0.56u
X335 a_n8659_n1230 a_n8537_n1530.t11 VSS.t89 VSS.t88 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X336 DEBUG.t67 a_n17351_68.t28 a_n15085_2072.t35 VSS.t272 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X337 VDD.t14 a_22388_3950.t5 a_22304_4398 VDD.t13 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X338 VDD.t271 PLL_DISABLE.t18 a_27899_438.t9 VDD.t270 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X339 a_24335_1611 a_22115_1610.t4 a_24090_1243 VSS.t120 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X340 PLL_CLK_OUT.t7 PLL_DISABLE.t19 a_24355_n1338.t15 VDD.t141 pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.33u
X341 a_23691_6933 a_n8537_n1530.t12 VSS.t321 VSS.t320 nfet_03v3 ad=0.26p pd=1.52u as=0.4p ps=1.8u w=1u l=0.33u
X342 a_22388_2038.t1 a_23508_2038 VDD.t73 VDD.t72 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X343 PLL_VCTRL.t19 PLL_FREERUN.t26 DEBUG.t13 VSS.t222 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X344 a_21394_11355.t9 a_21394_11355.t8 VDD.t174 VDD.t173 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X345 VDD.t143 PLL_DISABLE.t20 a_27899_438.t5 VDD.t142 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X346 a_1712_13773 a_5840_13333 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X347 a_24655_2486 a_24207_2486 VSS.t65 VSS.t64 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X348 a_24355_n1338.t16 PLL_DISABLE.t21 PLL_CLK_OUT.t8 VDD.t144 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X349 a_24090_1243 a_22527_1197 a_23455_1567 VSS.t66 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X350 a_21855_2486 a_21755_1082 VDD.t298 VDD.t297 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X351 a_22388_2038.t1 a_24655_2486 VDD.t99 VDD.t98 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X352 VDD.t193 a_21394_11355.t24 a_21506_13215.t3 VDD.t192 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X353 a_24355_n1338.t22 a_23423_n1258 VSS.t240 VSS.t239 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X354 DEBUG.t35 PLL_FREERUN.t27 a_n15085_2072.t5 VDD.t187 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X355 a_25369_6873 a_22388_2038.t3 VSS.t182 VSS.t181 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X356 a_22963_1518 a_24383_217 VDD.t93 VDD.t92 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X357 VSS.t261 a_n4208_n141.t5 a_14657_n1138 VSS.t260 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X358 a_24335_n301 a_22115_n302.t4 a_24090_n669 VSS.t108 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X359 a_22527_1197 a_22115_1610.t5 VDD.t358 VDD.t103 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X360 a_n2908_8493 a_1220_8933 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X361 DEBUG.t12 PLL_FREERUN.t28 PLL_VCTRL.t18 VSS.t336 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X362 a_1220_12453 a_5840_11573 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X363 VDD.t170 a_n8471_219.t9 a_14645_2840 VDD.t169 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X364 a_23427_n669 a_22115_n302.t5 a_23083_n301 VDD.t278 pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X365 a_25265_6933 a_26049_6873 a_26115_6933 VSS.t112 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X366 DEBUG.t71 a_n17351_68.t29 a_n15085_2072.t37 VSS.t314 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X367 a_23083_261 a_22963_217 a_22959_629 VDD.t59 pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X368 a_24090_n669 a_22527_n715 a_23455_n345 VSS.t58 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X369 a_23427_1243 a_22115_1610.t6 a_23083_1611 VDD.t102 pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X370 VDD.t71 a_23508_2038 a_22948_3950 VDD.t70 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X371 a_23508_2038 a_22304_4398 VDD.t24 VDD.t23 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X372 a_26795_7733 a_22941_7733.t5 a_25265_7733 VDD.t101 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X373 a_23691_6933 a_n8537_93.t9 a_23620_8319.t0 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X374 a_n2908_10253 a_1220_9813 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X375 a_21755_4907 a_21667_4951 VSS.t105 VSS.t104 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X376 a_5840_15093.t9 a_5840_7613.t0 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X377 a_25150_2082 a_24655_2486 VSS.t132 VSS.t131 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X378 a_22304_2486 a_22388_2038.t4 a_22324_2082 VSS.t269 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X379 PLL_VCTRL.t11 PLL_FREERUN.t29 DEBUG.t11 VSS.t337 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X380 a_n15085_2072.t4 PLL_FREERUN.t30 DEBUG.t34 VDD.t344 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X381 a_5840_15093.t9 a_5840_7613.t0 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X382 VDD.t161 a_22203_n358.t15 a_23423_n1258 VDD.t160 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X383 VSS.t263 a_n4208_n141.t6 a_3161_n1138 VSS.t262 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X384 a_27014_14933 a_27414_10401 VSS.t71 ppolyf_u r_width=0.8u r_length=22u
X385 a_24755_6933 a_24675_7463 VSS.t344 VSS.t343 nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.33u
X386 a_n15085_2072.t38 a_n17351_68.t30 DEBUG.t72 VSS.t315 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X387 a_1712_8493 a_5840_8933 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X388 VSS.t277 PLL_DISABLE.t22 a_27899_438.t6 VSS.t276 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X389 VSS.t215 a_22539_3430 a_22451_3522 VSS.t214 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X390 PLL_VCTRL.t10 PLL_FREERUN.t31 DEBUG.t10 VSS.t199 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X391 a_25675_1518 a_25587_1610 VDD.t319 VDD.t318 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X392 a_21394_11355.t7 a_21394_11355.t6 VDD.t255 VDD.t254 pfet_03v3 ad=1.456p pd=6.12u as=3.64p ps=12.5u w=5.6u l=0.56u
X393 VSS.t279 PLL_DISABLE.t23 a_27899_438.t7 VSS.t278 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X394 a_21891_6933 a_n8537_93.t10 a_n8537_n1530.t0 VSS.t46 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X395 VDD.t351 a_24675_7463 a_24755_6933 VDD.t350 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X396 a_21394_11355.t1 a_21506_13215.t11 a_24866_11400 VSS.t0 nfet_03v3 ad=1.456p pd=6.12u as=3.416p ps=12.42u w=5.6u l=0.56u
X397 VDD.t331 a_22864_4398 a_22388_3950.t0 VDD.t330 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X398 VDD.t253 a_21394_11355.t4 a_21394_11355.t5 VDD.t252 pfet_03v3 ad=3.64p pd=12.5u as=1.456p ps=6.12u w=5.6u l=0.56u
X399 VSS.t323 a_n8537_n1530.t13 a_26795_6933 VSS.t322 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X400 DEBUG.t73 a_n17351_68.t31 a_n15085_2072.t39 VSS.t316 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X401 DEBUG.t33 PLL_FREERUN.t32 a_n15085_2072.t3 VDD.t149 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X402 VSS.t209 a_22203_n358.t16 a_22115_253.t0 VSS.t207 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X403 PLL_CLK_OUT.t14 a_27899_438.t27 a_24355_n1338.t19 VSS.t221 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X404 a_n4208_n141.t1 a_n4208_n141.t0 VSS.t283 VSS.t282 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X405 a_24355_n1338.t49 a_27899_438.t28 PLL_CLK_OUT.t13 VSS.t349 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X406 DEBUG.t9 PLL_FREERUN.t33 PLL_VCTRL.t5 VSS.t200 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X407 VSS.t297 a_22987_3430 a_22899_3522 VSS.t296 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X408 a_22963_217 a_24383_n345 VSS.t11 VSS.t10 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X409 a_n8471_219.t1 a_n8537_93.t11 a_n8659_n1230 VSS.t116 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X410 a_24090_629 a_22527_574 a_23455_217 VSS.t58 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X411 VDD.t205 a_n8471_219.t10 a_6981_2840 VDD.t204 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X412 a_27899_438.t8 PLL_DISABLE.t24 VSS.t281 VSS.t280 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X413 a_5840_15093.t6 a_25369_6873 a_25265_6933 VSS.t291 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X414 VDD.t226 a_23423_n1258 a_24355_n1338.t30 VDD.t225 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X415 VSS.t238 a_23423_n1258 a_24355_n1338.t21 VSS.t237 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X416 a_1712_11133 a_5840_10693 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X417 a_n15085_2072.t2 PLL_FREERUN.t34 DEBUG.t32 VDD.t138 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X418 VDD.t88 PLL_DISABLE.t25 a_27899_438.t1 VDD.t87 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X419 a_n2908_14213 a_1220_13773 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
D2 VSS.t352 VDD.t53 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X420 a_n17351_68.t1 PLL_FREERUN.t35 VDD.t140 VDD.t139 pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.28u
X421 a_n15085_2072.t23 a_n17351_68.t32 DEBUG.t43 VSS.t158 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X422 VDD.t245 a_21394_11355.t2 a_21394_11355.t3 VDD.t244 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X423 VDD.t151 a_21394_11355.t25 a_n8537_n1530.t1 VDD.t150 pfet_03v3 ad=1.456p pd=5.78u as=0.5824p ps=2.76u w=2.24u l=0.56u
X424 a_23547_4907 a_23459_4951 VSS.t97 VSS.t96 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X425 a_25334_2082 a_22864_2486 a_25150_2082 VSS.t232 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X426 a_26115_6933 a_24675_7463 a_25265_7733 VDD.t349 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X427 VSS.t126 a_31479_1644 a_31391_1688 VSS.t125 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X428 VSS.t340 a_24383_1567 a_24335_1611 VSS.t339 nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X429 PLL_VCTRL.t4 PLL_FREERUN.t36 DEBUG.t8 VSS.t186 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X430 a_24355_n1338.t2 PLL_DISABLE.t26 PLL_CLK_OUT.t2 VDD.t89 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X431 VSS.t163 a_21643_3430 a_21555_3522 VSS.t162 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X432 a_11009_2840 a_7177_2840 a_10825_n1138 VSS.t80 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X433 a_24207_2486 a_22304_2486 VDD.t304 VDD.t303 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X434 a_n15085_2072.t48 VSS.t191 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X435 a_24706_3522 a_22304_2486 VSS.t303 VSS.t302 nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X436 VSS.t265 a_n4208_n141.t7 a_6993_n1138 VSS.t264 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X437 a_27899_438.t2 PLL_DISABLE.t27 VSS.t122 VSS.t121 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X438 a_23423_n1258 a_22203_n358.t17 VDD.t133 VDD.t132 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X439 DEBUG.t44 a_n17351_68.t33 a_n15085_2072.t24 VSS.t159 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X440 a_n2908_7613 a_1220_8053 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X441 VDD.t337 PLL_DISABLE.t28 a_27899_438.t10 VDD.t336 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X442 VSS.t9 a_24383_n345 a_24335_n301 VSS.t8 nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X443 a_22203_4907 a_22115_4951 VSS.t218 VSS.t217 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X444 a_27899_438.t11 PLL_DISABLE.t29 VSS.t329 VSS.t328 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X445 a_5840_15093.t9 VSS.t338 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X446 a_25675_n394 a_25587_n302 VDD.t288 VDD.t287 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X447 a_23995_4907 a_23907_4951 VSS.t180 VSS.t179 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X448 a_23423_n1258 a_22203_n358.t18 VDD.t135 VDD.t134 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X449 PLL_CLK_OUT.t12 a_27899_438.t29 a_24355_n1338.t50 VSS.t350 nfet_03v3 ad=0.26p pd=1.52u as=0.65p ps=3.3u w=1u l=0.33u
X450 a_24375_n669 a_22527_n715 a_24090_n669 VDD.t48 pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X451 a_22388_3950.t1 a_23508_2038 a_25334_3994 VSS.t81 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X452 a_24355_n1338.t51 a_27899_438.t30 PLL_CLK_OUT.t11 VSS.t351 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X453 a_24375_1243 a_22527_1197 a_24090_1243 VDD.t56 pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X454 PLL_CLK_OUT.t35 PLL_DISABLE.t30 a_24355_n1338.t48 VDD.t338 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X455 a_n8537_n1530.t2 a_21394_11355.t26 VDD.t153 VDD.t152 pfet_03v3 ad=0.5824p pd=2.76u as=0.5824p ps=2.76u w=2.24u l=0.56u
X456 a_21506_13215.t0 a_24866_11400 VSS.t1 VSS.t0 nfet_03v3 ad=1.456p pd=6.12u as=3.416p ps=12.42u w=5.6u l=0.56u
X457 a_24655_2486 a_24207_2486 VDD.t55 VDD.t54 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X458 a_21755_n830 a_21667_n786 VSS.t44 VSS.t43 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X459 a_n8659_n1230 a_n8537_n1530.t14 VSS.t5 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.33u
X460 a_n8659_n1230 a_n8537_93.t12 a_n8471_219.t1 VSS.t117 nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.33u
X461 a_24900_3522 a_22864_2486 a_24706_3522 VSS.t231 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X462 a_24355_n1338.t29 a_23423_n1258 VDD.t224 VDD.t223 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X463 PLL_CLK_OUT.t6 PLL_DISABLE.t31 a_24355_n1338.t14 VDD.t122 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X464 a_25369_6873 a_22388_2038.t5 VDD.t164 VDD.t163 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X465 a_26115_6933 a_24675_7463 a_25265_7733 VDD.t348 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X466 VDD.t222 a_23423_n1258 a_24355_n1338.t28 VDD.t221 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X467 a_5840_15093.t9 a_5840_7613.t0 cap_mim_2f0_m4m5_noshield c_width=11u c_length=11u
X468 a_27814_14933 VSS.t155 VSS.t154 ppolyf_u r_width=0.8u r_length=22u
X469 DEBUG.t45 a_n17351_68.t34 PLL_VCTRL.t21 VDD.t111 pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.33u
X470 a_25095_6933 a_n8537_n1530.t15 VSS.t7 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X471 a_22651_4907 a_22563_4951 VSS.t48 VSS.t47 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X472 a_22527_n715 a_22115_n302.t6 VSS.t197 VSS.t106 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X473 a_1712_7613 a_5840_8053 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X474 VSS.t174 PLL_DISABLE.t32 a_27899_438.t3 VSS.t173 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X475 a_25339_4907 a_25251_4951 VSS.t95 VSS.t94 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X476 DEBUG.t31 PLL_FREERUN.t37 a_n15085_2072.t1 VDD.t341 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X477 VSS.t228 a_n4208_n141.t8 a_10825_n1138 VSS.t227 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X478 DEBUG.t40 a_n17351_68.t35 a_n15085_2072.t21 VSS.t133 nfet_03v3 ad=0.65p pd=3.3u as=0.26p ps=1.52u w=1u l=0.33u
X479 a_n15085_2072.t22 a_n17351_68.t36 DEBUG.t41 VSS.t134 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X480 a_3345_2840 a_n487_2840 a_3161_n1138 VSS.t93 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X481 a_1712_10253 a_5840_9813 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
X482 a_n8537_93.t0 a_21394_11355.t27 VDD.t155 VDD.t154 pfet_03v3 ad=0.5824p pd=2.76u as=1.456p ps=5.78u w=2.24u l=0.56u
X483 a_23620_8319.t1 a_22941_7733.t6 a_23691_7733 VDD.t315 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X484 VDD.t137 a_22203_n358.t19 a_22115_n302.t1 VDD.t136 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X485 a_n2908_13333 a_1220_13333 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X486 VSS.t128 a_23435_3430 a_23347_3522 VSS.t127 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X487 a_27899_438.t4 PLL_DISABLE.t33 VSS.t176 VSS.t175 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X488 a_24355_n1338.t0 PLL_DISABLE.t34 PLL_CLK_OUT.t0 VDD.t62 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X489 a_n15085_2072.t49 VSS.t319 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X490 VSS.t290 a_25369_6873 a_26049_6873 VSS.t289 nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.33u
X491 a_24355_n1338.t20 a_23423_n1258 VSS.t236 VSS.t235 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X492 VSS.t51 a_21855_n1258 a_22203_n358.t0 VSS.t50 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X493 a_24090_n669 a_22115_n302.t7 a_23455_n345 VDD.t148 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X494 a_n15085_2072.t20 a_1220_14653 VSS.t17 ppolyf_u_1k r_width=1u r_length=20u
X495 VDD.t178 a_21394_11355.t28 a_n8537_93.t0 VDD.t177 pfet_03v3 ad=0.5824p pd=2.76u as=0.5824p ps=2.76u w=2.24u l=0.56u
X496 a_22884_3994 a_22304_4398 VSS.t32 VSS.t31 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X497 a_n15085_2072.t50 VSS.t190 cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
X498 a_24090_1243 a_22115_1610.t7 a_23455_1567 VDD.t86 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X499 a_21506_13215.t2 a_21394_11355.t29 VDD.t180 VDD.t179 pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X500 VSS.t75 PLL_DISABLE.t35 a_27899_438.t0 VSS.t74 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X501 a_24355_n1338.t6 a_27899_438.t31 PLL_CLK_OUT.t10 VSS.t156 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X502 a_22324_3994 a_21855_4398 VSS.t310 VSS.t309 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X503 PLL_CLK_OUT.t9 a_27899_438.t32 a_24355_n1338.t7 VSS.t157 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X504 DEBUG.t42 a_n17351_68.t37 PLL_VCTRL.t20 VDD.t105 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X505 VSS.t129 a_24383_217 a_24335_261 VSS.t8 nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X506 a_n8659_n1230 a_n8537_93.t13 a_n8471_219.t0 VSS.t330 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X507 VSS.t22 a_23883_3430 a_23795_3522 VSS.t21 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X508 PLL_CLK_OUT.t1 PLL_DISABLE.t36 a_24355_n1338.t1 VDD.t63 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X509 a_n17351_68.t0 PLL_FREERUN.t38 VSS.t333 VSS.t332 nfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
X510 a_5840_15093.t5 a_25369_6873 a_25265_6933 VSS.t288 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X511 PLL_VCTRL.t9 PLL_FREERUN.t39 DEBUG.t7 VSS.t334 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X512 a_n15085_2072.t25 a_n17351_68.t38 DEBUG.t46 VSS.t164 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X513 VSS.t26 a_27491_1710 a_21755_4018 VSS.t25 nfet_06v0 ad=0.151p pd=1.185u as=0.1261p ps=1.005u w=0.485u l=0.6u
X514 VDD.t207 a_n8471_219.t11 a_10813_2840 VDD.t206 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X515 a_n9701_6193 a_16431_6193 VSS.t183 ppolyf_u r_width=0.8u r_length=0.13m
X516 DEBUG.t30 PLL_FREERUN.t40 a_n15085_2072.t0 VDD.t237 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X517 a_24443_4907 a_24355_4951 VSS.t185 VSS.t184 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X518 a_n558_2704.t0 a_11009_2840 a_14645_2840 VDD.t147 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X519 PLL_VCTRL.t8 PLL_FREERUN.t41 DEBUG.t6 VSS.t253 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X520 a_25265_7733 a_24755_6933 a_5840_15093.t0 VDD.t125 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X521 PLL_VCTRL.t22 a_n17351_68.t39 DEBUG.t47 VDD.t117 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X522 a_1712_13773 a_5840_14213 VSS.t18 ppolyf_u_1k r_width=1u r_length=20u
D3 VSS.t187 PLL_DISABLE.t37 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X523 a_n8537_n1530.t3 a_n8537_93.t14 a_21891_6933 VSS.t331 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X524 DEBUG.t48 a_n17351_68.t40 PLL_VCTRL.t23 VDD.t118 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
X525 VSS.t208 a_22203_n358.t20 a_22115_n302.t0 VSS.t207 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X526 DEBUG.t61 a_n17351_68.t41 PLL_VCTRL.t30 VDD.t239 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.33u
R0 VSS.n3050 VSS.n158 108707
R1 VSS.n1651 VSS.n1078 71567.2
R2 VSS.n3050 VSS.n159 63487.1
R3 VSS.n1604 VSS.n1092 57292.9
R4 VSS.n1653 VSS.t109 44684.9
R5 VSS.n1558 VSS.n1557 41487.9
R6 VSS.n1588 VSS.n1587 41443.1
R7 VSS.n1653 VSS.n1072 40731.1
R8 VSS.n1441 VSS.n1440 38820.7
R9 VSS.n1654 VSS.n1653 38116.5
R10 VSS.n1652 VSS.n1651 17415.5
R11 VSS.t27 VSS.n1092 13315.1
R12 VSS.n1652 VSS.n1077 13283.7
R13 VSS.n1605 VSS.n1604 12117.8
R14 VSS.n138 VSS.n18 12018.2
R15 VSS.n838 VSS.n158 11767.2
R16 VSS.n873 VSS.n838 11262.4
R17 VSS.n3481 VSS.n3480 10496.9
R18 VSS.n1587 VSS.n1558 8427.59
R19 VSS.n2302 VSS.n556 8157.71
R20 VSS.n466 VSS.n435 8157.71
R21 VSS.n2569 VSS.n313 8157.71
R22 VSS.n2747 VSS.n353 8157.71
R23 VSS.n1606 VSS.n1605 8040.81
R24 VSS.n1653 VSS.n1652 7822.41
R25 VSS.n3101 VSS.n99 7592.86
R26 VSS.n1392 VSS.n1108 7347.33
R27 VSS.n2216 VSS.n555 7312.98
R28 VSS.n2960 VSS.n203 7297.55
R29 VSS.t150 VSS.n3467 6174.11
R30 VSS.n2961 VSS.n2960 5958.33
R31 VSS.n140 VSS.n139 4966.24
R32 VSS.n203 VSS.n202 4966.24
R33 VSS.n3476 VSS.n3475 4888.01
R34 VSS.n1557 VSS.n1556 4674.55
R35 VSS.n1603 VSS.n1405 4606.25
R36 VSS.n1440 VSS.n1078 4034.48
R37 VSS.n1622 VSS.n1092 3728.12
R38 VSS.n142 VSS.n138 3373.39
R39 VSS.n3467 VSS.n18 2712.26
R40 VSS.n139 VSS.n81 2681.51
R41 VSS.n9 VSS.t148 2585.85
R42 VSS.n3476 VSS.n9 2574.44
R43 VSS.n789 VSS.n18 2530.6
R44 VSS.t183 VSS.n81 2437.5
R45 VSS.n3475 VSS.n10 2409.43
R46 VSS.n3453 VSS.n34 2232.27
R47 VSS.n34 VSS.n9 2232.27
R48 VSS.n3158 VSS.n37 1975.11
R49 VSS.n3480 VSS.n6 1861.31
R50 VSS.n1603 VSS.t241 1799.8
R51 VSS.n1624 VSS.n1623 1756.25
R52 VSS.n1606 VSS.n1404 1755.41
R53 VSS.t203 VSS.t299 1662.1
R54 VSS.t29 VSS.n1405 1565.64
R55 VSS.n3478 VSS.n6 1540.41
R56 VSS.t43 VSS.t207 1513.7
R57 VSS.n3158 VSS.t183 1503.17
R58 VSS.n1623 VSS.n1622 1493.75
R59 VSS.n139 VSS.n117 1460.46
R60 VSS.t36 VSS.t10 1439.5
R61 VSS.n3453 VSS.t271 1421.85
R62 VSS.n1588 VSS.n1441 1412.07
R63 VSS.t131 VSS.t171 1406.11
R64 VSS.t177 VSS.t90 1394.98
R65 VSS.t106 VSS.t151 1365.3
R66 VSS.n194 VSS.t282 1362.36
R67 VSS.n1623 VSS.t181 1298.52
R68 VSS.n1586 VSS.t43 1261.42
R69 VSS.t306 VSS.t19 1250.29
R70 VSS.t10 VSS.n1585 1246.58
R71 VSS.n1559 VSS.t29 1231.74
R72 VSS.t67 VSS.t308 1202.05
R73 VSS.t14 VSS.t59 1202.05
R74 VSS.n1389 VSS.n1108 1192.59
R75 VSS.n40 VSS.t198 1191.86
R76 VSS.n947 VSS.n615 1186.87
R77 VSS.n947 VSS.n946 1171.01
R78 VSS.t40 VSS.t12 1157.53
R79 VSS.n1389 VSS.n1388 1146.55
R80 VSS.n1402 VSS.n1108 1125.34
R81 VSS.n1604 VSS.n1603 1122.18
R82 VSS.n1123 VSS.t23 1113.01
R83 VSS.n1439 VSS.t299 1113.01
R84 VSS.t84 VSS.n1124 1109.3
R85 VSS.t296 VSS.t326 1101.88
R86 VSS.t83 VSS.t15 1101.88
R87 VSS.t239 VSS.t201 1044.49
R88 VSS.t311 VSS.t56 1044.49
R89 VSS.n1390 VSS.n1389 1029.84
R90 VSS.t8 VSS.t36 994.293
R91 VSS.n3453 VSS.n3452 982.053
R92 VSS.t332 VSS.n10 982.053
R93 VSS.t38 VSS.t82 960.903
R94 VSS.n1513 VSS.t212 949.024
R95 VSS.n2360 VSS.t260 949.024
R96 VSS.n2394 VSS.t227 949.024
R97 VSS.n2627 VSS.t264 949.024
R98 VSS.n2661 VSS.t262 949.024
R99 VSS.n255 VSS.t210 949.024
R100 VSS.n793 VSS.n789 908.319
R101 VSS.n1440 VSS.n589 904.097
R102 VSS.n3467 VSS.t133 899.178
R103 VSS.t52 VSS.t229 889.111
R104 VSS.n1513 VSS.t226 873.673
R105 VSS.n2360 VSS.t196 873.673
R106 VSS.n2394 VSS.t80 873.673
R107 VSS.n2627 VSS.t92 873.673
R108 VSS.n2661 VSS.t93 873.673
R109 VSS.n255 VSS.t266 873.673
R110 VSS.n2216 VSS.n589 868.476
R111 VSS.n1125 VSS.t162 845.89
R112 VSS.n1122 VSS.n1121 831.051
R113 VSS.t58 VSS.t108 831.051
R114 VSS.t12 VSS.t58 831.051
R115 VSS.t207 VSS.t106 831.051
R116 VSS.n1390 VSS.n1090 807.538
R117 VSS.n3463 VSS.t99 782.889
R118 VSS.n14 VSS.t192 769.885
R119 VSS.t325 VSS.t81 756.85
R120 VSS.t231 VSS.t33 756.85
R121 VSS.n1405 VSS.n1092 753.125
R122 VSS.n1120 VSS.n1119 749.429
R123 VSS.n1589 VSS.n1588 728.482
R124 VSS.t302 VSS.t231 719.75
R125 VSS.n1125 VSS.n1078 719.75
R126 VSS.n1441 VSS.n1439 719.75
R127 VSS.n1587 VSS.n1586 719.75
R128 VSS.t49 VSS.t214 708.62
R129 VSS.t214 VSS.t31 686.359
R130 VSS.t21 VSS.t34 682.649
R131 VSS.t31 VSS.t153 682.649
R132 VSS.t309 VSS.t49 682.649
R133 VSS.t66 VSS.n1419 682.649
R134 VSS.t269 VSS.t69 682.649
R135 VSS.n3466 VSS.n19 657.931
R136 VSS.t232 VSS.t341 649.259
R137 VSS.n1411 VSS.t311 647.41
R138 VSS.n850 VSS.n849 643.222
R139 VSS.t64 VSS.t339 638.129
R140 VSS.n1423 VSS.t232 626.999
R141 VSS.t339 VSS.t120 623.288
R142 VSS.t108 VSS.t8 623.288
R143 VSS.t59 VSS.t40 623.288
R144 VSS.t151 VSS.t14 623.288
R145 VSS.t125 VSS.t285 588.216
R146 VSS.n3026 VSS.n3025 583.484
R147 VSS.n3025 VSS.n3024 583.484
R148 VSS.n3024 VSS.n2998 583.484
R149 VSS.n3018 VSS.n2998 583.484
R150 VSS.n3018 VSS.n3017 583.484
R151 VSS.n3017 VSS.n3016 583.484
R152 VSS.n3016 VSS.n3002 583.484
R153 VSS.n3010 VSS.n3002 583.484
R154 VSS.n3010 VSS.n3009 583.484
R155 VSS.n3009 VSS.n3008 583.484
R156 VSS.n3008 VSS.n5 583.484
R157 VSS.n3481 VSS.n5 583.484
R158 VSS.n3026 VSS.n2997 583.271
R159 VSS.t216 VSS.t118 567.638
R160 VSS.n3101 VSS.n117 564.85
R161 VSS.t326 VSS.t127 560.217
R162 VSS.n847 VSS.n21 552.693
R163 VSS.t72 VSS.n1120 549.087
R164 VSS.t77 VSS.t324 549.087
R165 VSS.t34 VSS.n1123 549.087
R166 VSS.n1555 VSS.n1446 534.539
R167 VSS.n1549 VSS.n1548 534.539
R168 VSS.n1548 VSS.n1547 534.539
R169 VSS.n1547 VSS.n1507 534.539
R170 VSS.n1541 VSS.n1507 534.539
R171 VSS.n1541 VSS.n1540 534.539
R172 VSS.n1540 VSS.n1539 534.539
R173 VSS.n1539 VSS.n1511 534.539
R174 VSS.n1532 VSS.n1511 534.539
R175 VSS.n1532 VSS.n1531 534.539
R176 VSS.n1531 VSS.n1530 534.539
R177 VSS.n1530 VSS.n1516 534.539
R178 VSS.n1524 VSS.n1516 534.539
R179 VSS.n1524 VSS.n1523 534.539
R180 VSS.n1523 VSS.n1522 534.539
R181 VSS.n1522 VSS.n533 534.539
R182 VSS.n2340 VSS.n533 534.539
R183 VSS.n2347 VSS.n2346 534.539
R184 VSS.n2348 VSS.n2347 534.539
R185 VSS.n2348 VSS.n524 534.539
R186 VSS.n2354 VSS.n524 534.539
R187 VSS.n2355 VSS.n2354 534.539
R188 VSS.n2356 VSS.n2355 534.539
R189 VSS.n2356 VSS.n520 534.539
R190 VSS.n2364 VSS.n520 534.539
R191 VSS.n2365 VSS.n2364 534.539
R192 VSS.n2366 VSS.n2365 534.539
R193 VSS.n2366 VSS.n516 534.539
R194 VSS.n2372 VSS.n516 534.539
R195 VSS.n2373 VSS.n2372 534.539
R196 VSS.n2374 VSS.n2373 534.539
R197 VSS.n2374 VSS.n512 534.539
R198 VSS.n2380 VSS.n512 534.539
R199 VSS.n2381 VSS.n2380 534.539
R200 VSS.n2382 VSS.n2381 534.539
R201 VSS.n2436 VSS.n497 534.539
R202 VSS.n2430 VSS.n497 534.539
R203 VSS.n2430 VSS.n2429 534.539
R204 VSS.n2429 VSS.n2428 534.539
R205 VSS.n2428 VSS.n2388 534.539
R206 VSS.n2422 VSS.n2388 534.539
R207 VSS.n2422 VSS.n2421 534.539
R208 VSS.n2421 VSS.n2420 534.539
R209 VSS.n2420 VSS.n2392 534.539
R210 VSS.n2413 VSS.n2392 534.539
R211 VSS.n2413 VSS.n2412 534.539
R212 VSS.n2412 VSS.n2411 534.539
R213 VSS.n2411 VSS.n2397 534.539
R214 VSS.n2405 VSS.n2397 534.539
R215 VSS.n2405 VSS.n2404 534.539
R216 VSS.n2404 VSS.n2403 534.539
R217 VSS.n2403 VSS.n413 534.539
R218 VSS.n2607 VSS.n413 534.539
R219 VSS.n2614 VSS.n2613 534.539
R220 VSS.n2615 VSS.n2614 534.539
R221 VSS.n2615 VSS.n404 534.539
R222 VSS.n2621 VSS.n404 534.539
R223 VSS.n2622 VSS.n2621 534.539
R224 VSS.n2623 VSS.n2622 534.539
R225 VSS.n2623 VSS.n400 534.539
R226 VSS.n2631 VSS.n400 534.539
R227 VSS.n2632 VSS.n2631 534.539
R228 VSS.n2633 VSS.n2632 534.539
R229 VSS.n2633 VSS.n396 534.539
R230 VSS.n2639 VSS.n396 534.539
R231 VSS.n2640 VSS.n2639 534.539
R232 VSS.n2641 VSS.n2640 534.539
R233 VSS.n2641 VSS.n392 534.539
R234 VSS.n2647 VSS.n392 534.539
R235 VSS.n2648 VSS.n2647 534.539
R236 VSS.n2649 VSS.n2648 534.539
R237 VSS.n2708 VSS.n379 534.539
R238 VSS.n2702 VSS.n379 534.539
R239 VSS.n2702 VSS.n2701 534.539
R240 VSS.n2701 VSS.n2700 534.539
R241 VSS.n2700 VSS.n2655 534.539
R242 VSS.n2694 VSS.n2655 534.539
R243 VSS.n2694 VSS.n2693 534.539
R244 VSS.n2693 VSS.n2692 534.539
R245 VSS.n2692 VSS.n2659 534.539
R246 VSS.n2685 VSS.n2659 534.539
R247 VSS.n2685 VSS.n2684 534.539
R248 VSS.n2684 VSS.n2683 534.539
R249 VSS.n2683 VSS.n2664 534.539
R250 VSS.n2677 VSS.n2664 534.539
R251 VSS.n2677 VSS.n2676 534.539
R252 VSS.n2676 VSS.n2675 534.539
R253 VSS.n2675 VSS.n2668 534.539
R254 VSS.n2668 VSS.n267 534.539
R255 VSS.n2881 VSS.n262 534.539
R256 VSS.n2887 VSS.n262 534.539
R257 VSS.n2888 VSS.n2887 534.539
R258 VSS.n2889 VSS.n2888 534.539
R259 VSS.n2889 VSS.n258 534.539
R260 VSS.n2895 VSS.n258 534.539
R261 VSS.n2896 VSS.n2895 534.539
R262 VSS.n2897 VSS.n2896 534.539
R263 VSS.n2897 VSS.n253 534.539
R264 VSS.n2904 VSS.n253 534.539
R265 VSS.n2905 VSS.n2904 534.539
R266 VSS.n2906 VSS.n2905 534.539
R267 VSS.n2906 VSS.n249 534.539
R268 VSS.n2912 VSS.n249 534.539
R269 VSS.n2913 VSS.n2912 534.539
R270 VSS.n2914 VSS.n2913 534.539
R271 VSS.n2914 VSS.n243 534.539
R272 VSS.n2937 VSS.n2936 534.539
R273 VSS.n2936 VSS.n2935 534.539
R274 VSS.n2935 VSS.n2928 534.539
R275 VSS.t116 VSS.t117 519.268
R276 VSS.t330 VSS.t116 519.268
R277 VSS.t99 VSS.t330 519.268
R278 VSS.t142 VSS.t4 510.158
R279 VSS.t88 VSS.t142 510.158
R280 VSS.t192 VSS.t88 510.158
R281 VSS.n1549 VSS.n1506 494.45
R282 VSS.t123 VSS.t233 486.017
R283 VSS.t104 VSS.n1644 484.224
R284 VSS.t241 VSS.t243 483.401
R285 VSS.t243 VSS.t247 483.401
R286 VSS.t247 VSS.t235 483.401
R287 VSS.t235 VSS.t245 483.401
R288 VSS.t245 VSS.t249 483.401
R289 VSS.t249 VSS.t237 483.401
R290 VSS.t237 VSS.t239 483.401
R291 VSS.t229 VSS.t205 483.401
R292 VSS.t54 VSS.t52 483.401
R293 VSS.t50 VSS.t54 483.401
R294 VSS.t56 VSS.t50 483.401
R295 VSS.t183 VSS.n80 444.149
R296 VSS.n3451 VSS.n37 435.764
R297 VSS.n1124 VSS.t21 430.365
R298 VSS.t304 VSS.t66 430.365
R299 VSS.n1557 VSS.n1411 418.659
R300 VSS.n1359 VSS.n1355 416.675
R301 VSS.n1284 VSS.n1267 403.765
R302 VSS.n1284 VSS.n1283 403.765
R303 VSS.n1283 VSS.n1282 403.765
R304 VSS.n1282 VSS.n1268 403.765
R305 VSS.n1276 VSS.n1268 403.765
R306 VSS.n1276 VSS.n1275 403.765
R307 VSS.n1275 VSS.n1076 403.765
R308 VSS.t120 VSS.t304 400.685
R309 VSS.n1645 VSS.t144 394.5
R310 VSS.n2214 VSS.n2213 388.524
R311 VSS.n2217 VSS.n583 388.524
R312 VSS.n2223 VSS.n583 388.524
R313 VSS.n2224 VSS.n2223 388.524
R314 VSS.n2225 VSS.n2224 388.524
R315 VSS.n2225 VSS.n579 388.524
R316 VSS.n2231 VSS.n579 388.524
R317 VSS.n2232 VSS.n2231 388.524
R318 VSS.n2233 VSS.n2232 388.524
R319 VSS.n2233 VSS.n575 388.524
R320 VSS.n2239 VSS.n575 388.524
R321 VSS.n2240 VSS.n2239 388.524
R322 VSS.n2241 VSS.n2240 388.524
R323 VSS.n2241 VSS.n571 388.524
R324 VSS.n2247 VSS.n571 388.524
R325 VSS.n2248 VSS.n2247 388.524
R326 VSS.n2249 VSS.n2248 388.524
R327 VSS.n2301 VSS.n557 388.524
R328 VSS.n2295 VSS.n557 388.524
R329 VSS.n2295 VSS.n2294 388.524
R330 VSS.n2294 VSS.n2293 388.524
R331 VSS.n2293 VSS.n2255 388.524
R332 VSS.n2287 VSS.n2255 388.524
R333 VSS.n2287 VSS.n2286 388.524
R334 VSS.n2286 VSS.n2285 388.524
R335 VSS.n2285 VSS.n2259 388.524
R336 VSS.n2279 VSS.n2259 388.524
R337 VSS.n2279 VSS.n2278 388.524
R338 VSS.n2278 VSS.n2277 388.524
R339 VSS.n2277 VSS.n2263 388.524
R340 VSS.n2271 VSS.n2263 388.524
R341 VSS.n2271 VSS.n2270 388.524
R342 VSS.n2270 VSS.n2269 388.524
R343 VSS.n2269 VSS.n472 388.524
R344 VSS.n2471 VSS.n472 388.524
R345 VSS.n2478 VSS.n2477 388.524
R346 VSS.n2479 VSS.n2478 388.524
R347 VSS.n2479 VSS.n462 388.524
R348 VSS.n2485 VSS.n462 388.524
R349 VSS.n2486 VSS.n2485 388.524
R350 VSS.n2487 VSS.n2486 388.524
R351 VSS.n2487 VSS.n458 388.524
R352 VSS.n2493 VSS.n458 388.524
R353 VSS.n2494 VSS.n2493 388.524
R354 VSS.n2495 VSS.n2494 388.524
R355 VSS.n2495 VSS.n454 388.524
R356 VSS.n2501 VSS.n454 388.524
R357 VSS.n2502 VSS.n2501 388.524
R358 VSS.n2503 VSS.n2502 388.524
R359 VSS.n2503 VSS.n450 388.524
R360 VSS.n2509 VSS.n450 388.524
R361 VSS.n2510 VSS.n2509 388.524
R362 VSS.n2511 VSS.n2510 388.524
R363 VSS.n2568 VSS.n436 388.524
R364 VSS.n2562 VSS.n436 388.524
R365 VSS.n2562 VSS.n2561 388.524
R366 VSS.n2561 VSS.n2560 388.524
R367 VSS.n2560 VSS.n2517 388.524
R368 VSS.n2554 VSS.n2517 388.524
R369 VSS.n2554 VSS.n2553 388.524
R370 VSS.n2553 VSS.n2552 388.524
R371 VSS.n2552 VSS.n2521 388.524
R372 VSS.n2546 VSS.n2521 388.524
R373 VSS.n2546 VSS.n2545 388.524
R374 VSS.n2545 VSS.n2544 388.524
R375 VSS.n2544 VSS.n2525 388.524
R376 VSS.n2538 VSS.n2525 388.524
R377 VSS.n2538 VSS.n2537 388.524
R378 VSS.n2537 VSS.n2536 388.524
R379 VSS.n2536 VSS.n2529 388.524
R380 VSS.n2529 VSS.n355 388.524
R381 VSS.n2749 VSS.n2748 388.524
R382 VSS.n2749 VSS.n307 388.524
R383 VSS.n2755 VSS.n307 388.524
R384 VSS.n2756 VSS.n2755 388.524
R385 VSS.n2757 VSS.n2756 388.524
R386 VSS.n2757 VSS.n303 388.524
R387 VSS.n2763 VSS.n303 388.524
R388 VSS.n2764 VSS.n2763 388.524
R389 VSS.n2765 VSS.n2764 388.524
R390 VSS.n2765 VSS.n299 388.524
R391 VSS.n2771 VSS.n299 388.524
R392 VSS.n2772 VSS.n2771 388.524
R393 VSS.n2773 VSS.n2772 388.524
R394 VSS.n2773 VSS.n295 388.524
R395 VSS.n2780 VSS.n295 388.524
R396 VSS.n2781 VSS.n2780 388.524
R397 VSS.n2782 VSS.n2781 388.524
R398 VSS.n2782 VSS.n285 388.524
R399 VSS.n2831 VSS.n2830 388.524
R400 VSS.n2830 VSS.n2829 388.524
R401 VSS.n2829 VSS.n2788 388.524
R402 VSS.n2823 VSS.n2788 388.524
R403 VSS.n2823 VSS.n2822 388.524
R404 VSS.n2822 VSS.n2821 388.524
R405 VSS.n2821 VSS.n2792 388.524
R406 VSS.n2815 VSS.n2792 388.524
R407 VSS.n2815 VSS.n2814 388.524
R408 VSS.n2814 VSS.n2813 388.524
R409 VSS.n2813 VSS.n2796 388.524
R410 VSS.n2807 VSS.n2796 388.524
R411 VSS.n2807 VSS.n2806 388.524
R412 VSS.n2806 VSS.n2805 388.524
R413 VSS.n2805 VSS.n2800 388.524
R414 VSS.n2800 VSS.n118 388.524
R415 VSS.n3093 VSS.n3092 388.524
R416 VSS.n3092 VSS.n3091 388.524
R417 VSS.n3091 VSS.n130 388.524
R418 VSS.t222 VSS.t150 387.993
R419 VSS.t223 VSS.t222 387.993
R420 VSS.t199 VSS.t223 387.993
R421 VSS.t318 VSS.t199 387.993
R422 VSS.t273 VSS.t318 387.993
R423 VSS.t268 VSS.t273 387.993
R424 VSS.t149 VSS.t268 387.993
R425 VSS.t336 VSS.t149 387.993
R426 VSS.t225 VSS.t336 387.993
R427 VSS.t200 VSS.t253 387.993
R428 VSS.t253 VSS.t275 387.993
R429 VSS.t275 VSS.t334 387.993
R430 VSS.t337 VSS.t274 387.993
R431 VSS.t317 VSS.t337 387.993
R432 VSS.t186 VSS.t317 387.993
R433 VSS.t259 VSS.t186 387.993
R434 VSS.t148 VSS.t259 387.993
R435 VSS.n1359 VSS.n614 384.562
R436 VSS.n2944 VSS.n243 379.524
R437 VSS.n1607 VSS.n1107 375.974
R438 VSS.n1461 VSS.n590 372.921
R439 VSS.n1476 VSS.n1461 372.921
R440 VSS.n1477 VSS.n1476 372.921
R441 VSS.n1479 VSS.n1477 372.921
R442 VSS.n1479 VSS.n1478 372.921
R443 VSS.n1478 VSS.n1442 372.921
R444 VSS.n1456 VSS.n1443 372.921
R445 VSS.n1490 VSS.n1456 372.921
R446 VSS.n1491 VSS.n1490 372.921
R447 VSS.n1492 VSS.n1491 372.921
R448 VSS.n1492 VSS.n1451 372.921
R449 VSS.n1505 VSS.n1451 372.921
R450 VSS.n2928 VSS.n238 366.161
R451 VSS.n202 VSS.n133 364.974
R452 VSS.t86 VSS.n1638 361.745
R453 VSS.t171 VSS.t64 356.164
R454 VSS.n873 VSS.n872 354.031
R455 VSS.n872 VSS.n871 354.031
R456 VSS.n871 VSS.n839 354.031
R457 VSS.n865 VSS.n839 354.031
R458 VSS.n865 VSS.n864 354.031
R459 VSS.n1558 VSS.n1442 346.817
R460 VSS.n864 VSS.n17 341.639
R461 VSS.n1392 VSS.n1391 336.921
R462 VSS.n2216 VSS.n2215 336.074
R463 VSS.n1625 VSS.n1090 334.796
R464 VSS.n3429 VSS.n3158 332.938
R465 VSS.n1556 VSS.n1555 331.414
R466 VSS.n2937 VSS.n244 331.414
R467 VSS.n1602 VSS.t205 328.022
R468 VSS.n1506 VSS.n1505 324.442
R469 VSS.n3101 VSS.n118 316.647
R470 VSS.n224 VSS.n223 316.457
R471 VSS.n230 VSS.n210 316.457
R472 VSS.n231 VSS.n230 316.457
R473 VSS.n232 VSS.n231 316.457
R474 VSS.n232 VSS.n204 316.457
R475 VSS.n2959 VSS.n205 316.457
R476 VSS.n2953 VSS.n205 316.457
R477 VSS.n2953 VSS.n2952 316.457
R478 VSS.n2952 VSS.n2951 316.457
R479 VSS.n2945 VSS.n242 316.457
R480 VSS.t25 VSS.t27 315.973
R481 VSS.n889 VSS.n793 310.856
R482 VSS.n1304 VSS.n1303 308.411
R483 VSS.n1303 VSS.n1302 308.411
R484 VSS.n1302 VSS.n1294 308.411
R485 VSS.n1296 VSS.n1294 308.411
R486 VSS.n1296 VSS.n1075 308.411
R487 VSS.n1654 VSS.n1075 308.411
R488 VSS.n2346 VSS.n528 307.361
R489 VSS.n2437 VSS.n2436 307.361
R490 VSS.n2613 VSS.n408 307.361
R491 VSS.n2709 VSS.n2708 307.361
R492 VSS.n2881 VSS.n2880 307.361
R493 VSS.n1589 VSS.n591 306.935
R494 VSS.t96 VSS.t194 306.202
R495 VSS.n2963 VSS.n2962 302.748
R496 VSS.n2963 VSS.n197 302.748
R497 VSS.n2970 VSS.n197 302.748
R498 VSS.n2971 VSS.n2970 302.748
R499 VSS.n2972 VSS.n2971 302.748
R500 VSS.n2972 VSS.n192 302.748
R501 VSS.n2978 VSS.n192 302.748
R502 VSS.n2979 VSS.n2978 302.748
R503 VSS.n2980 VSS.n2979 302.748
R504 VSS.n2980 VSS.n188 302.748
R505 VSS.n2986 VSS.n188 302.748
R506 VSS.n2987 VSS.n2986 302.748
R507 VSS.n2988 VSS.n2987 302.748
R508 VSS.n3040 VSS.n171 302.748
R509 VSS.n3034 VSS.n171 302.748
R510 VSS.n3034 VSS.n3033 302.748
R511 VSS.n3033 VSS.n3032 302.748
R512 VSS.n3032 VSS.n159 296.693
R513 VSS.t153 VSS.t296 293.094
R514 VSS.t274 VSS.n6 289.853
R515 VSS.n3467 VSS.n3466 288.923
R516 VSS.n2340 VSS.n2339 288.651
R517 VSS.n2382 VSS.n496 288.651
R518 VSS.n2607 VSS.n2606 288.651
R519 VSS.n2649 VSS.n378 288.651
R520 VSS.n2879 VSS.n267 288.651
R521 VSS.n2943 VSS.n244 288.651
R522 VSS.n3469 VSS.n15 286.461
R523 VSS.n3460 VSS.n20 286.447
R524 VSS.n1121 VSS.t72 281.964
R525 VSS.n139 VSS.n138 277.757
R526 VSS.n3057 VSS.n152 277.659
R527 VSS.n3051 VSS.n152 277.659
R528 VSS.n3049 VSS.n3048 277.659
R529 VSS.n3048 VSS.n160 277.659
R530 VSS.t134 VSS.t133 275.425
R531 VSS.t168 VSS.t134 275.425
R532 VSS.t315 VSS.t168 275.425
R533 VSS.t335 VSS.t315 275.425
R534 VSS.t158 VSS.t335 275.425
R535 VSS.t257 VSS.t158 275.425
R536 VSS.t164 VSS.t257 275.425
R537 VSS.t272 VSS.t164 275.425
R538 VSS.t267 VSS.t272 275.425
R539 VSS.t284 VSS.t170 275.425
R540 VSS.t270 VSS.t284 275.425
R541 VSS.t258 VSS.t270 275.425
R542 VSS.t314 VSS.t258 275.425
R543 VSS.t169 VSS.t314 275.425
R544 VSS.t316 VSS.t169 275.425
R545 VSS.t224 VSS.t316 275.425
R546 VSS.t159 VSS.t224 275.425
R547 VSS.t271 VSS.t159 275.425
R548 VSS.n2945 VSS.n2944 275.317
R549 VSS.n2960 VSS.n2959 273.735
R550 VSS.n1267 VSS.n1077 272.236
R551 VSS.t90 VSS.t309 270.834
R552 VSS.n2304 VSS.n548 270.495
R553 VSS.n2310 VSS.n548 270.495
R554 VSS.n2311 VSS.n2310 270.495
R555 VSS.n2312 VSS.n2311 270.495
R556 VSS.n2312 VSS.n544 270.495
R557 VSS.n2318 VSS.n544 270.495
R558 VSS.n2319 VSS.n2318 270.495
R559 VSS.n2320 VSS.n2319 270.495
R560 VSS.n2320 VSS.n540 270.495
R561 VSS.n2326 VSS.n540 270.495
R562 VSS.n2327 VSS.n2326 270.495
R563 VSS.n2329 VSS.n2327 270.495
R564 VSS.n2329 VSS.n2328 270.495
R565 VSS.n2463 VSS.n2462 270.495
R566 VSS.n2462 VSS.n2461 270.495
R567 VSS.n2461 VSS.n484 270.495
R568 VSS.n2455 VSS.n484 270.495
R569 VSS.n2455 VSS.n2454 270.495
R570 VSS.n2454 VSS.n2453 270.495
R571 VSS.n2453 VSS.n488 270.495
R572 VSS.n2447 VSS.n488 270.495
R573 VSS.n2447 VSS.n2446 270.495
R574 VSS.n2446 VSS.n2445 270.495
R575 VSS.n2445 VSS.n492 270.495
R576 VSS.n2439 VSS.n492 270.495
R577 VSS.n2439 VSS.n2438 270.495
R578 VSS.n2571 VSS.n428 270.495
R579 VSS.n2577 VSS.n428 270.495
R580 VSS.n2578 VSS.n2577 270.495
R581 VSS.n2579 VSS.n2578 270.495
R582 VSS.n2579 VSS.n424 270.495
R583 VSS.n2585 VSS.n424 270.495
R584 VSS.n2586 VSS.n2585 270.495
R585 VSS.n2587 VSS.n2586 270.495
R586 VSS.n2587 VSS.n420 270.495
R587 VSS.n2593 VSS.n420 270.495
R588 VSS.n2594 VSS.n2593 270.495
R589 VSS.n2596 VSS.n2594 270.495
R590 VSS.n2596 VSS.n2595 270.495
R591 VSS.n2734 VSS.n354 270.495
R592 VSS.n2734 VSS.n2733 270.495
R593 VSS.n2733 VSS.n2732 270.495
R594 VSS.n2732 VSS.n365 270.495
R595 VSS.n2726 VSS.n365 270.495
R596 VSS.n2726 VSS.n2725 270.495
R597 VSS.n2725 VSS.n2724 270.495
R598 VSS.n2724 VSS.n370 270.495
R599 VSS.n2718 VSS.n370 270.495
R600 VSS.n2718 VSS.n2717 270.495
R601 VSS.n2717 VSS.n2716 270.495
R602 VSS.n2716 VSS.n374 270.495
R603 VSS.n2710 VSS.n374 270.495
R604 VSS.n2843 VSS.n281 270.495
R605 VSS.n2849 VSS.n281 270.495
R606 VSS.n2850 VSS.n2849 270.495
R607 VSS.n2851 VSS.n2850 270.495
R608 VSS.n2851 VSS.n277 270.495
R609 VSS.n2857 VSS.n277 270.495
R610 VSS.n2858 VSS.n2857 270.495
R611 VSS.n2859 VSS.n2858 270.495
R612 VSS.n2859 VSS.n273 270.495
R613 VSS.n2865 VSS.n273 270.495
R614 VSS.n2866 VSS.n2865 270.495
R615 VSS.n2867 VSS.n2866 270.495
R616 VSS.n2867 VSS.n266 270.495
R617 VSS.t162 VSS.t177 267.123
R618 VSS.t15 VSS.t181 267.123
R619 VSS.n2213 VSS.n591 264.197
R620 VSS.n3093 VSS.n129 264.197
R621 VSS.n3058 VSS.n3057 263.776
R622 VSS.t81 VSS.n1122 255.994
R623 VSS.t343 VSS.t184 254.93
R624 VSS.n1613 VSS.n1102 253.106
R625 VSS.n1611 VSS.n1103 253.106
R626 VSS.n1406 VSS.n1107 253.106
R627 VSS.n3469 VSS.n16 253.106
R628 VSS.n3460 VSS.n24 253.106
R629 VSS.n3100 VSS.n119 252.541
R630 VSS.n1391 VSS.n1093 249.606
R631 VSS.n1613 VSS.n1094 249.606
R632 VSS.n1611 VSS.n1104 249.606
R633 VSS.n3458 VSS.n25 249.606
R634 VSS.n3458 VSS.n26 249.606
R635 VSS.n3452 VSS.n3451 245.012
R636 VSS.t102 VSS.t47 243.536
R637 VSS.n19 VSS.n17 242.852
R638 VSS.n202 VSS.n130 242.827
R639 VSS.t294 VSS.t291 242.113
R640 VSS.t288 VSS.t140 242.113
R641 VSS.t140 VSS.t6 242.113
R642 VSS.t345 VSS.t343 242.113
R643 VSS.t139 VSS.t45 242.113
R644 VSS.t194 VSS.t141 242.113
R645 VSS.t138 VSS.t102 242.113
R646 VSS.t46 VSS.t331 242.113
R647 VSS.t331 VSS.t100 242.113
R648 VSS.n3050 VSS.n3049 240.175
R649 VSS.t167 VSS.t255 239.8
R650 VSS.t286 VSS.t156 239.8
R651 VSS.t351 VSS.t220 239.8
R652 VSS.t165 VSS.t254 239.8
R653 VSS.t166 VSS.t256 239.8
R654 VSS.t157 VSS.t349 239.8
R655 VSS.t276 VSS.t219 238.391
R656 VSS.n2302 VSS.n2301 237
R657 VSS.n2477 VSS.n466 237
R658 VSS.n2569 VSS.n2568 237
R659 VSS.n2748 VSS.n2747 237
R660 VSS.n2831 VSS.n99 237
R661 VSS.n2328 VSS.n528 235.332
R662 VSS.n2438 VSS.n2437 235.332
R663 VSS.n2595 VSS.n408 235.332
R664 VSS.n2710 VSS.n2709 235.332
R665 VSS.n2880 VSS.n266 235.332
R666 VSS.t63 VSS.t295 232.143
R667 VSS.t136 VSS.t280 229.927
R668 VSS.n3474 VSS.n7 226.763
R669 VSS.t350 VSS.t25 221.464
R670 VSS.n1355 VSS.n1352 207.988
R671 VSS.n1304 VSS.n1077 207.945
R672 VSS.n3076 VSS.n3075 207.668
R673 VSS.n3075 VSS.n3074 207.668
R674 VSS.n3074 VSS.n143 207.668
R675 VSS.n3068 VSS.n143 207.668
R676 VSS.n3068 VSS.n3067 207.668
R677 VSS.n3067 VSS.n3066 207.668
R678 VSS.n3066 VSS.n147 207.668
R679 VSS.n3060 VSS.n147 207.668
R680 VSS.n3060 VSS.n3059 207.668
R681 VSS.n887 VSS.n794 207.668
R682 VSS.n881 VSS.n794 207.668
R683 VSS.n881 VSS.n880 207.668
R684 VSS.n880 VSS.n879 207.668
R685 VSS.n1401 VSS.t286 201.714
R686 VSS.t82 VSS.t123 196.632
R687 VSS.t60 VSS.t167 196.072
R688 VSS.n1402 VSS.t125 194.661
R689 VSS.n3468 VSS.t225 193.996
R690 VSS.n3468 VSS.t200 193.996
R691 VSS.n879 VSS.n158 191.054
R692 VSS.t295 VSS.t94 189.417
R693 VSS.n3041 VSS.n3040 187.704
R694 VSS.n2249 VSS.n552 186.492
R695 VSS.n2471 VSS.n2470 186.492
R696 VSS.n2511 VSS.n432 186.492
R697 VSS.n2745 VSS.n355 186.492
R698 VSS.n2841 VSS.n285 186.492
R699 VSS.n129 VSS.n128 186.492
R700 VSS.n1625 VSS.t289 176.279
R701 VSS.t173 VSS.t137 173.504
R702 VSS.n2951 VSS.n238 172.469
R703 VSS.t33 VSS.t77 170.662
R704 VSS.t221 VSS.t328 165.04
R705 VSS.n224 VSS.n203 164.558
R706 VSS.n1119 VSS.t115 163.782
R707 VSS.t121 VSS.t135 162.219
R708 VSS.n1161 VSS.t68 161.487
R709 VSS.n1098 VSS.t287 159.398
R710 VSS.n2961 VSS.n201 158.944
R711 VSS.t201 VSS.n1602 155.379
R712 VSS.n2944 VSS.n2943 155.017
R713 VSS.t251 VSS.t138 152.388
R714 VSS.n210 VSS.n203 151.899
R715 VSS.n1645 VSS.t47 150.964
R716 VSS.t278 VSS.t221 150.934
R717 VSS.t217 VSS.t46 149.541
R718 VSS.n1419 VSS.t38 148.403
R719 VSS.n1384 VSS.t154 148.343
R720 VSS.t42 VSS.n1153 147.215
R721 VSS.n1404 VSS.n1402 145.553
R722 VSS.t146 VSS.t350 145.292
R723 VSS.t19 VSS.t269 144.692
R724 VSS.n242 VSS.n238 143.988
R725 VSS.n1639 VSS.t320 143.844
R726 VSS.n2962 VSS.n2961 143.805
R727 VSS.t137 VSS.t175 142.47
R728 VSS.t71 VSS.n1381 141.207
R729 VSS.t347 VSS.t345 140.995
R730 VSS.t187 VSS.t157 139.649
R731 VSS.n1637 VSS.t184 139.571
R732 VSS.t45 VSS.t179 138.147
R733 VSS.n3459 VSS.t267 137.713
R734 VSS.n3459 VSS.t170 137.713
R735 VSS.t233 VSS.t67 137.273
R736 VSS.n128 VSS.n119 135.983
R737 VSS.n3482 VSS.n4 135.464
R738 VSS.t324 VSS.t325 133.562
R739 VSS.n141 VSS.n140 131.869
R740 VSS.n1423 VSS.t83 129.852
R741 VSS.n142 VSS.n141 129.792
R742 VSS.n889 VSS.n888 124.343
R743 VSS.t115 VSS.n1118 123.904
R744 VSS.n1607 VSS.n1103 122.868
R745 VSS.n3474 VSS.n11 122.868
R746 VSS.n33 VSS.n24 122.868
R747 VSS.n33 VSS.n16 122.868
R748 VSS.t127 VSS.t84 122.433
R749 VSS.n1612 VSS.t135 119.9
R750 VSS.n1118 VSS.t294 118.209
R751 VSS.t23 VSS.t302 115.011
R752 VSS.t118 VSS.t306 115.011
R753 VSS.t289 VSS.t292 108.186
R754 VSS.t292 VSS.t322 108.186
R755 VSS.t322 VSS.t98 108.186
R756 VSS.t114 VSS.t112 108.186
R757 VSS.t113 VSS.t114 108.186
R758 VSS.t179 VSS.t86 103.966
R759 VSS.n16 VSS.n7 103.895
R760 VSS.n36 VSS.n24 103.895
R761 VSS.n36 VSS.n11 103.895
R762 VSS.t6 VSS.t347 101.118
R763 VSS.t287 VSS.t187 100.153
R764 VSS.n140 VSS.n133 99.9337
R765 VSS.n1375 VSS.n1162 99.1454
R766 VSS.n1369 VSS.n1162 99.1454
R767 VSS.n1369 VSS.n1368 99.1454
R768 VSS.n1368 VSS.n1367 99.1454
R769 VSS.n1362 VSS.n1361 99.1454
R770 VSS.n1351 VSS.n1222 99.1454
R771 VSS.n1345 VSS.n1222 99.1454
R772 VSS.n1290 VSS.n1228 99.1454
R773 VSS.n1639 VSS.t139 98.2696
R774 VSS.t334 VSS.n6 98.1395
R775 VSS.t175 VSS.t166 97.3312
R776 VSS.n238 VSS.n201 95.3661
R777 VSS.n905 VSS.n904 94.601
R778 VSS.n904 VSS.n903 94.601
R779 VSS.n903 VSS.n785 94.601
R780 VSS.n897 VSS.n785 94.601
R781 VSS.t349 VSS.t146 94.51
R782 VSS.t144 VSS.t217 92.5728
R783 VSS.t141 VSS.t251 89.7244
R784 VSS.t156 VSS.t278 88.8677
R785 VSS.n2988 VSS.n167 87.7974
R786 VSS.n1093 VSS.n1091 87.1213
R787 VSS.n1601 VSS.n1406 86.2755
R788 VSS.t74 VSS.t136 86.0465
R789 VSS.n1601 VSS.n1407 82.7755
R790 VSS.n1361 VSS.n1360 82.6213
R791 VSS.t256 VSS.n1098 80.4041
R792 VSS.n1624 VSS.t112 79.5482
R793 VSS.n1392 VSS.n1102 77.9216
R794 VSS.n3076 VSS.n142 77.8759
R795 VSS.n888 VSS.n151 77.8759
R796 VSS.t219 VSS.t121 77.583
R797 VSS.n3041 VSS.n167 75.6875
R798 VSS.t328 VSS.t351 74.7618
R799 VSS.n1406 VSS.n1104 74.1422
R800 VSS.n3101 VSS.n3100 71.8774
R801 VSS.n1345 VSS.n1344 69.8526
R802 VSS.t254 VSS.t173 66.2982
R803 VSS.n1375 VSS.n1161 65.346
R804 VSS.n3467 VSS.n17 64.4305
R805 VSS.n2154 VSS.n614 63.438
R806 VSS.n888 VSS.n887 63.3392
R807 VSS.n1641 VSS.n1640 62.7954
R808 VSS.n1652 VSS.n1061 60.9861
R809 VSS.n167 VSS.n160 59.6972
R810 VSS.t308 VSS.t216 55.6512
R811 VSS.n1660 VSS.n1659 54.8952
R812 VSS.n1376 VSS.n1159 53.1452
R813 VSS.n2172 VSS.n587 53.0314
R814 VSS.n2165 VSS.n588 53.0314
R815 VSS.n2165 VSS.n2164 53.0314
R816 VSS.n2164 VSS.n2163 53.0314
R817 VSS.n2163 VSS.n608 53.0314
R818 VSS.n2157 VSS.n608 53.0314
R819 VSS.n2157 VSS.n2156 53.0314
R820 VSS.n2149 VSS.n2148 53.0314
R821 VSS.n2148 VSS.n2147 53.0314
R822 VSS.n2147 VSS.n1762 53.0314
R823 VSS.n2141 VSS.n1762 53.0314
R824 VSS.n2141 VSS.n2140 53.0314
R825 VSS.n2140 VSS.n2139 53.0314
R826 VSS.n2139 VSS.n1767 53.0314
R827 VSS.n2133 VSS.n1767 53.0314
R828 VSS.n2133 VSS.n2132 53.0314
R829 VSS.n1815 VSS.n554 53.0314
R830 VSS.n2124 VSS.n1815 53.0314
R831 VSS.n2124 VSS.n2123 53.0314
R832 VSS.n2123 VSS.n2122 53.0314
R833 VSS.n2122 VSS.n1816 53.0314
R834 VSS.n2116 VSS.n1816 53.0314
R835 VSS.n2116 VSS.n2115 53.0314
R836 VSS.n2115 VSS.n2114 53.0314
R837 VSS.n2114 VSS.n1820 53.0314
R838 VSS.n2108 VSS.n1820 53.0314
R839 VSS.n2108 VSS.n2107 53.0314
R840 VSS.n2107 VSS.n2106 53.0314
R841 VSS.n2106 VSS.n1824 53.0314
R842 VSS.n2100 VSS.n1824 53.0314
R843 VSS.n2100 VSS.n2099 53.0314
R844 VSS.n2099 VSS.n2098 53.0314
R845 VSS.n2098 VSS.n1828 53.0314
R846 VSS.n2092 VSS.n1828 53.0314
R847 VSS.n2050 VSS.n2049 53.0314
R848 VSS.n2049 VSS.n2048 53.0314
R849 VSS.n2048 VSS.n1833 53.0314
R850 VSS.n2042 VSS.n1833 53.0314
R851 VSS.n2042 VSS.n2041 53.0314
R852 VSS.n2041 VSS.n2040 53.0314
R853 VSS.n2040 VSS.n1838 53.0314
R854 VSS.n2034 VSS.n1838 53.0314
R855 VSS.n2034 VSS.n2033 53.0314
R856 VSS.n2033 VSS.n2032 53.0314
R857 VSS.n2032 VSS.n1842 53.0314
R858 VSS.n2026 VSS.n1842 53.0314
R859 VSS.n2026 VSS.n2025 53.0314
R860 VSS.n2025 VSS.n2024 53.0314
R861 VSS.n2024 VSS.n1846 53.0314
R862 VSS.n2018 VSS.n1846 53.0314
R863 VSS.n2018 VSS.n2017 53.0314
R864 VSS.n2017 VSS.n2016 53.0314
R865 VSS.n2009 VSS.n434 53.0314
R866 VSS.n2009 VSS.n2008 53.0314
R867 VSS.n2008 VSS.n2007 53.0314
R868 VSS.n2007 VSS.n1894 53.0314
R869 VSS.n2001 VSS.n1894 53.0314
R870 VSS.n2001 VSS.n2000 53.0314
R871 VSS.n2000 VSS.n1999 53.0314
R872 VSS.n1999 VSS.n1899 53.0314
R873 VSS.n1993 VSS.n1899 53.0314
R874 VSS.n1993 VSS.n1992 53.0314
R875 VSS.n1992 VSS.n1991 53.0314
R876 VSS.n1991 VSS.n1903 53.0314
R877 VSS.n1985 VSS.n1903 53.0314
R878 VSS.n1985 VSS.n1984 53.0314
R879 VSS.n1984 VSS.n1983 53.0314
R880 VSS.n1983 VSS.n1907 53.0314
R881 VSS.n1977 VSS.n1907 53.0314
R882 VSS.n1977 VSS.n1976 53.0314
R883 VSS.n1954 VSS.n312 53.0314
R884 VSS.n1968 VSS.n1954 53.0314
R885 VSS.n1968 VSS.n1967 53.0314
R886 VSS.n1967 VSS.n1966 53.0314
R887 VSS.n1966 VSS.n1955 53.0314
R888 VSS.n1960 VSS.n1955 53.0314
R889 VSS.n1959 VSS.n79 53.0314
R890 VSS.n3151 VSS.n88 53.0314
R891 VSS.n3151 VSS.n3150 53.0314
R892 VSS.n3150 VSS.n3149 53.0314
R893 VSS.n3149 VSS.n89 53.0314
R894 VSS.n3143 VSS.n89 53.0314
R895 VSS.n3143 VSS.n3142 53.0314
R896 VSS.n3142 VSS.n3141 53.0314
R897 VSS.n3141 VSS.n93 53.0314
R898 VSS.n3134 VSS.n3133 53.0314
R899 VSS.n3133 VSS.n3132 53.0314
R900 VSS.n3132 VSS.n100 53.0314
R901 VSS.n3126 VSS.n100 53.0314
R902 VSS.n3126 VSS.n3125 53.0314
R903 VSS.n3125 VSS.n3124 53.0314
R904 VSS.n3124 VSS.n104 53.0314
R905 VSS.n3118 VSS.n104 53.0314
R906 VSS.n3118 VSS.n3117 53.0314
R907 VSS.n3117 VSS.n3116 53.0314
R908 VSS.n3110 VSS.n111 53.0314
R909 VSS.n3110 VSS.n3109 53.0314
R910 VSS.n3109 VSS.n3108 53.0314
R911 VSS.n3108 VSS.n112 53.0314
R912 VSS.n3102 VSS.n112 53.0314
R913 VSS.n743 VSS.n116 53.0314
R914 VSS.n750 VSS.n749 53.0314
R915 VSS.n751 VSS.n750 53.0314
R916 VSS.n751 VSS.n70 53.0314
R917 VSS.n1374 VSS.n1163 52.7768
R918 VSS.n88 VSS.n82 52.7663
R919 VSS.t94 VSS.t288 52.6955
R920 VSS.n1652 VSS.n1076 52.0005
R921 VSS.n3058 VSS.n151 51.9174
R922 VSS.n905 VSS.n80 51.0848
R923 VSS.n1352 VSS.n1083 50.2036
R924 VSS.n2216 VSS.n587 49.8496
R925 VSS.n1644 VSS.t109 49.8471
R926 VSS.n3059 VSS.n3058 47.7641
R927 VSS.n2217 VSS.n2216 46.6233
R928 VSS.n3102 VSS.n3101 46.4026
R929 VSS.t285 VSS.t60 43.7288
R930 VSS.n1621 VSS.n1093 43.1088
R931 VSS.n2960 VSS.n204 42.722
R932 VSS.t183 VSS.n79 42.4252
R933 VSS.n1248 VSS.n1218 40.5598
R934 VSS.n1506 VSS.n1446 40.091
R935 VSS.n1960 VSS.t18 40.0388
R936 VSS.n2210 VSS.n593 39.3485
R937 VSS.n1448 VSS.n593 39.3305
R938 VSS.n31 VSS.n10 38.8471
R939 VSS.n2156 VSS.n2155 38.4479
R940 VSS.t255 VSS.n1401 38.0864
R941 VSS.n3452 VSS.t332 37.9805
R942 VSS.n3051 VSS.n3050 37.4845
R943 VSS.n1311 VSS.n1310 37.0268
R944 VSS.n3116 VSS.t17 36.857
R945 VSS.n1343 VSS.n1226 36.6584
R946 VSS.n1690 VSS.n1061 36.0615
R947 VSS.n1403 VSS.n1102 35.6452
R948 VSS.n1403 VSS.n1103 35.6452
R949 VSS.n3454 VSS.n32 35.6452
R950 VSS.n3454 VSS.n24 35.6452
R951 VSS.n32 VSS.n31 35.6452
R952 VSS.n31 VSS.n11 35.6452
R953 VSS.n1119 VSS.t113 35.0015
R954 VSS.n1612 VSS.t74 33.8547
R955 VSS.t2 VSS.n1210 33.4243
R956 VSS.n1251 VSS.t0 33.4243
R957 VSS.t341 VSS.t131 33.3909
R958 VSS.n2173 VSS.n2172 32.8797
R959 VSS.n749 VSS.n700 32.8797
R960 VSS.n1638 VSS.n1637 32.7569
R961 VSS.n1290 VSS.n1077 32.2977
R962 VSS.n1367 VSS.n1210 31.9222
R963 VSS.n1691 VSS.n1059 30.5794
R964 VSS.n3479 VSS.n4 30.2813
R965 VSS.n2209 VSS.n595 29.7905
R966 VSS.n2210 VSS.n2209 29.7725
R967 VSS.n1585 VSS.n1559 29.6809
R968 VSS.n1344 VSS.n1228 29.2933
R969 VSS.n2302 VSS.n554 29.1675
R970 VSS.n2050 VSS.n466 29.1675
R971 VSS.n2569 VSS.n434 29.1675
R972 VSS.n2747 VSS.n312 29.1675
R973 VSS.n3134 VSS.n99 29.1675
R974 VSS.t98 VSS.n1624 28.6377
R975 VSS.n2132 VSS.n553 28.6372
R976 VSS.n2092 VSS.n2091 28.6372
R977 VSS.n2016 VSS.n433 28.6372
R978 VSS.n1976 VSS.n311 28.6372
R979 VSS.n743 VSS.n700 28.6372
R980 VSS.n1688 VSS.n1070 28.3689
R981 VSS.n1684 VSS.n1683 28.3689
R982 VSS.n1680 VSS.n1679 28.3689
R983 VSS.n1676 VSS.n1675 28.3689
R984 VSS.n1672 VSS.n1671 28.3689
R985 VSS.n1668 VSS.n1667 28.3689
R986 VSS.n1664 VSS.n1663 28.3689
R987 VSS.n1201 VSS.n1199 28.0005
R988 VSS.n1199 VSS.n1198 28.0005
R989 VSS.n1195 VSS.n1194 28.0005
R990 VSS.n1192 VSS.n1168 28.0005
R991 VSS.n1188 VSS.n1186 28.0005
R992 VSS.n1184 VSS.n1170 28.0005
R993 VSS.n1180 VSS.n1178 28.0005
R994 VSS.n1176 VSS.n1173 28.0005
R995 VSS.n1343 VSS.n1237 28.0005
R996 VSS.n1339 VSS.n1338 28.0005
R997 VSS.n1335 VSS.n1334 28.0005
R998 VSS.n1331 VSS.n1330 28.0005
R999 VSS.n1327 VSS.n1326 28.0005
R1000 VSS.n1323 VSS.n1322 28.0005
R1001 VSS.n1319 VSS.n1318 28.0005
R1002 VSS.n1315 VSS.n1314 28.0005
R1003 VSS.n3478 VSS.n3477 27.5094
R1004 VSS.n1252 VSS.n1241 26.6645
R1005 VSS.n1558 VSS.n1443 26.1049
R1006 VSS.n1104 VSS.n1094 24.7922
R1007 VSS.n1374 VSS.n1164 24.3163
R1008 VSS.n1370 VSS.n1164 24.3163
R1009 VSS.n1370 VSS.n1206 24.3163
R1010 VSS.n1366 VSS.n1206 24.3163
R1011 VSS.n1363 VSS.n1211 24.3163
R1012 VSS.n1363 VSS.n1217 24.3163
R1013 VSS.n1350 VSS.n1217 24.3163
R1014 VSS.n1350 VSS.n1223 24.3163
R1015 VSS.n1346 VSS.n1223 24.3163
R1016 VSS.n1289 VSS.n1262 24.3163
R1017 VSS.n1289 VSS.n1263 24.3163
R1018 VSS.n1285 VSS.n1263 24.3163
R1019 VSS.n1285 VSS.n1266 24.3163
R1020 VSS.n1281 VSS.n1266 24.3163
R1021 VSS.n1281 VSS.n1269 24.3163
R1022 VSS.n1277 VSS.n1269 24.3163
R1023 VSS.n1277 VSS.n1274 24.3163
R1024 VSS.n1274 VSS.n1273 24.3163
R1025 VSS.n1273 VSS.n1059 24.3163
R1026 VSS.n1376 VSS.n1160 24.3163
R1027 VSS.n1207 VSS.n1160 24.3163
R1028 VSS.n1208 VSS.n1207 24.3163
R1029 VSS.n1209 VSS.n1208 24.3163
R1030 VSS.n1253 VSS.n1209 24.3163
R1031 VSS.n1253 VSS.n1219 24.3163
R1032 VSS.n1220 VSS.n1219 24.3163
R1033 VSS.n1221 VSS.n1220 24.3163
R1034 VSS.n1258 VSS.n1221 24.3163
R1035 VSS.n1258 VSS.n1227 24.3163
R1036 VSS.n1309 VSS.n1291 24.3163
R1037 VSS.n1305 VSS.n1291 24.3163
R1038 VSS.n1305 VSS.n1293 24.3163
R1039 VSS.n1301 VSS.n1293 24.3163
R1040 VSS.n1301 VSS.n1295 24.3163
R1041 VSS.n1297 VSS.n1295 24.3163
R1042 VSS.n1297 VSS.n1074 24.3163
R1043 VSS.n1655 VSS.n1074 24.3163
R1044 VSS.n1655 VSS.n1072 24.3163
R1045 VSS.n1659 VSS.n1072 24.3163
R1046 VSS.n1691 VSS.n1060 24.2242
R1047 VSS.n1649 VSS.t110 24.116
R1048 VSS.n2339 VSS.n528 24.0548
R1049 VSS.n2437 VSS.n496 24.0548
R1050 VSS.n2606 VSS.n408 24.0548
R1051 VSS.n2709 VSS.n378 24.0548
R1052 VSS.n2880 VSS.n2879 24.0548
R1053 VSS.n1637 VSS.n1636 23.9005
R1054 VSS.n1646 VSS.n1645 23.9005
R1055 VSS.n2302 VSS.n555 23.7479
R1056 VSS.n556 VSS.n466 23.7479
R1057 VSS.n2569 VSS.n435 23.7479
R1058 VSS.n2747 VSS.n313 23.7479
R1059 VSS.n353 VSS.n99 23.7479
R1060 VSS.n1648 VSS.t101 22.3205
R1061 VSS.n1647 VSS.t145 22.3205
R1062 VSS.n1080 VSS.t103 22.3205
R1063 VSS.n1635 VSS.t87 22.3205
R1064 VSS.n1632 VSS.t344 22.3205
R1065 VSS.n1627 VSS.t290 22.3205
R1066 VSS.n1062 VSS.n603 21.2129
R1067 VSS.n2173 VSS.n603 20.6826
R1068 VSS.n1634 VSS.n1633 19.8005
R1069 VSS.n1631 VSS.n1630 19.8005
R1070 VSS.n1629 VSS.n1628 19.8005
R1071 VSS.n897 VSS.n18 18.9206
R1072 VSS.n564 VSS.n563 18.4216
R1073 VSS.n2305 VSS.n551 18.4216
R1074 VSS.n2305 VSS.n549 18.4216
R1075 VSS.n2309 VSS.n549 18.4216
R1076 VSS.n2309 VSS.n547 18.4216
R1077 VSS.n2313 VSS.n547 18.4216
R1078 VSS.n2313 VSS.n545 18.4216
R1079 VSS.n2317 VSS.n545 18.4216
R1080 VSS.n2317 VSS.n543 18.4216
R1081 VSS.n2321 VSS.n543 18.4216
R1082 VSS.n2321 VSS.n541 18.4216
R1083 VSS.n2325 VSS.n541 18.4216
R1084 VSS.n2325 VSS.n539 18.4216
R1085 VSS.n2330 VSS.n539 18.4216
R1086 VSS.n2330 VSS.n537 18.4216
R1087 VSS.n2337 VSS.n537 18.4216
R1088 VSS.n2333 VSS.n536 18.4216
R1089 VSS.n2468 VSS.n480 18.4216
R1090 VSS.n2464 VSS.n479 18.4216
R1091 VSS.n2464 VSS.n483 18.4216
R1092 VSS.n2460 VSS.n483 18.4216
R1093 VSS.n2460 VSS.n485 18.4216
R1094 VSS.n2456 VSS.n485 18.4216
R1095 VSS.n2456 VSS.n487 18.4216
R1096 VSS.n2452 VSS.n487 18.4216
R1097 VSS.n2452 VSS.n489 18.4216
R1098 VSS.n2448 VSS.n489 18.4216
R1099 VSS.n2448 VSS.n491 18.4216
R1100 VSS.n2444 VSS.n491 18.4216
R1101 VSS.n2444 VSS.n493 18.4216
R1102 VSS.n2440 VSS.n493 18.4216
R1103 VSS.n2440 VSS.n495 18.4216
R1104 VSS.n503 VSS.n495 18.4216
R1105 VSS.n506 VSS.n505 18.4216
R1106 VSS.n443 VSS.n442 18.4216
R1107 VSS.n2572 VSS.n431 18.4216
R1108 VSS.n2572 VSS.n429 18.4216
R1109 VSS.n2576 VSS.n429 18.4216
R1110 VSS.n2576 VSS.n427 18.4216
R1111 VSS.n2580 VSS.n427 18.4216
R1112 VSS.n2580 VSS.n425 18.4216
R1113 VSS.n2584 VSS.n425 18.4216
R1114 VSS.n2584 VSS.n423 18.4216
R1115 VSS.n2588 VSS.n423 18.4216
R1116 VSS.n2588 VSS.n421 18.4216
R1117 VSS.n2592 VSS.n421 18.4216
R1118 VSS.n2592 VSS.n419 18.4216
R1119 VSS.n2597 VSS.n419 18.4216
R1120 VSS.n2597 VSS.n417 18.4216
R1121 VSS.n2604 VSS.n417 18.4216
R1122 VSS.n2600 VSS.n416 18.4216
R1123 VSS.n2739 VSS.n359 18.4216
R1124 VSS.n2737 VSS.n2736 18.4216
R1125 VSS.n2736 VSS.n2735 18.4216
R1126 VSS.n2735 VSS.n363 18.4216
R1127 VSS.n2731 VSS.n363 18.4216
R1128 VSS.n2731 VSS.n366 18.4216
R1129 VSS.n2727 VSS.n366 18.4216
R1130 VSS.n2727 VSS.n369 18.4216
R1131 VSS.n2723 VSS.n369 18.4216
R1132 VSS.n2723 VSS.n371 18.4216
R1133 VSS.n2719 VSS.n371 18.4216
R1134 VSS.n2719 VSS.n373 18.4216
R1135 VSS.n2715 VSS.n373 18.4216
R1136 VSS.n2715 VSS.n375 18.4216
R1137 VSS.n2711 VSS.n375 18.4216
R1138 VSS.n2711 VSS.n377 18.4216
R1139 VSS.n386 VSS.n385 18.4216
R1140 VSS.n2835 VSS.n289 18.4216
R1141 VSS.n2844 VSS.n284 18.4216
R1142 VSS.n2844 VSS.n282 18.4216
R1143 VSS.n2848 VSS.n282 18.4216
R1144 VSS.n2848 VSS.n280 18.4216
R1145 VSS.n2852 VSS.n280 18.4216
R1146 VSS.n2852 VSS.n278 18.4216
R1147 VSS.n2856 VSS.n278 18.4216
R1148 VSS.n2856 VSS.n276 18.4216
R1149 VSS.n2860 VSS.n276 18.4216
R1150 VSS.n2860 VSS.n274 18.4216
R1151 VSS.n2864 VSS.n274 18.4216
R1152 VSS.n2864 VSS.n272 18.4216
R1153 VSS.n2868 VSS.n272 18.4216
R1154 VSS.n2868 VSS.n270 18.4216
R1155 VSS.n2877 VSS.n270 18.4216
R1156 VSS.n2873 VSS.n269 18.4216
R1157 VSS.n828 VSS.n827 18.4216
R1158 VSS.n824 VSS.n823 18.4216
R1159 VSS.n821 VSS.n818 18.4216
R1160 VSS.n3056 VSS.n153 18.4216
R1161 VSS.n3056 VSS.n154 18.4216
R1162 VSS.n3052 VSS.n154 18.4216
R1163 VSS.n3052 VSS.n157 18.4216
R1164 VSS.n3047 VSS.n157 18.4216
R1165 VSS.n3047 VSS.n161 18.4216
R1166 VSS.n3043 VSS.n161 18.4216
R1167 VSS.n174 VSS.n166 18.4216
R1168 VSS.n178 VSS.n177 18.4216
R1169 VSS.n182 VSS.n181 18.4216
R1170 VSS.n1554 VSS.n1447 18.4216
R1171 VSS.n1550 VSS.n1447 18.4216
R1172 VSS.n1550 VSS.n1450 18.4216
R1173 VSS.n1546 VSS.n1450 18.4216
R1174 VSS.n1546 VSS.n1508 18.4216
R1175 VSS.n1542 VSS.n1508 18.4216
R1176 VSS.n1542 VSS.n1510 18.4216
R1177 VSS.n1538 VSS.n1510 18.4216
R1178 VSS.n1538 VSS.n1512 18.4216
R1179 VSS.n1533 VSS.n1512 18.4216
R1180 VSS.n1533 VSS.n1515 18.4216
R1181 VSS.n1529 VSS.n1515 18.4216
R1182 VSS.n1529 VSS.n1517 18.4216
R1183 VSS.n1525 VSS.n1517 18.4216
R1184 VSS.n1525 VSS.n1519 18.4216
R1185 VSS.n1521 VSS.n1519 18.4216
R1186 VSS.n1521 VSS.n532 18.4216
R1187 VSS.n2341 VSS.n532 18.4216
R1188 VSS.n2345 VSS.n527 18.4216
R1189 VSS.n2349 VSS.n527 18.4216
R1190 VSS.n2349 VSS.n525 18.4216
R1191 VSS.n2353 VSS.n525 18.4216
R1192 VSS.n2353 VSS.n523 18.4216
R1193 VSS.n2357 VSS.n523 18.4216
R1194 VSS.n2357 VSS.n521 18.4216
R1195 VSS.n2363 VSS.n521 18.4216
R1196 VSS.n2363 VSS.n519 18.4216
R1197 VSS.n2367 VSS.n519 18.4216
R1198 VSS.n2367 VSS.n517 18.4216
R1199 VSS.n2371 VSS.n517 18.4216
R1200 VSS.n2371 VSS.n515 18.4216
R1201 VSS.n2375 VSS.n515 18.4216
R1202 VSS.n2375 VSS.n513 18.4216
R1203 VSS.n2379 VSS.n513 18.4216
R1204 VSS.n2379 VSS.n511 18.4216
R1205 VSS.n2383 VSS.n511 18.4216
R1206 VSS.n2435 VSS.n499 18.4216
R1207 VSS.n2431 VSS.n499 18.4216
R1208 VSS.n2431 VSS.n2387 18.4216
R1209 VSS.n2427 VSS.n2387 18.4216
R1210 VSS.n2427 VSS.n2389 18.4216
R1211 VSS.n2423 VSS.n2389 18.4216
R1212 VSS.n2423 VSS.n2391 18.4216
R1213 VSS.n2419 VSS.n2391 18.4216
R1214 VSS.n2419 VSS.n2393 18.4216
R1215 VSS.n2414 VSS.n2393 18.4216
R1216 VSS.n2414 VSS.n2396 18.4216
R1217 VSS.n2410 VSS.n2396 18.4216
R1218 VSS.n2410 VSS.n2398 18.4216
R1219 VSS.n2406 VSS.n2398 18.4216
R1220 VSS.n2406 VSS.n2400 18.4216
R1221 VSS.n2402 VSS.n2400 18.4216
R1222 VSS.n2402 VSS.n412 18.4216
R1223 VSS.n2608 VSS.n412 18.4216
R1224 VSS.n2612 VSS.n407 18.4216
R1225 VSS.n2616 VSS.n407 18.4216
R1226 VSS.n2616 VSS.n405 18.4216
R1227 VSS.n2620 VSS.n405 18.4216
R1228 VSS.n2620 VSS.n403 18.4216
R1229 VSS.n2624 VSS.n403 18.4216
R1230 VSS.n2624 VSS.n401 18.4216
R1231 VSS.n2630 VSS.n401 18.4216
R1232 VSS.n2630 VSS.n399 18.4216
R1233 VSS.n2634 VSS.n399 18.4216
R1234 VSS.n2634 VSS.n397 18.4216
R1235 VSS.n2638 VSS.n397 18.4216
R1236 VSS.n2638 VSS.n395 18.4216
R1237 VSS.n2642 VSS.n395 18.4216
R1238 VSS.n2642 VSS.n393 18.4216
R1239 VSS.n2646 VSS.n393 18.4216
R1240 VSS.n2646 VSS.n391 18.4216
R1241 VSS.n2650 VSS.n391 18.4216
R1242 VSS.n2707 VSS.n381 18.4216
R1243 VSS.n2703 VSS.n381 18.4216
R1244 VSS.n2703 VSS.n2654 18.4216
R1245 VSS.n2699 VSS.n2654 18.4216
R1246 VSS.n2699 VSS.n2656 18.4216
R1247 VSS.n2695 VSS.n2656 18.4216
R1248 VSS.n2695 VSS.n2658 18.4216
R1249 VSS.n2691 VSS.n2658 18.4216
R1250 VSS.n2691 VSS.n2660 18.4216
R1251 VSS.n2686 VSS.n2660 18.4216
R1252 VSS.n2686 VSS.n2663 18.4216
R1253 VSS.n2682 VSS.n2663 18.4216
R1254 VSS.n2682 VSS.n2665 18.4216
R1255 VSS.n2678 VSS.n2665 18.4216
R1256 VSS.n2678 VSS.n2667 18.4216
R1257 VSS.n2674 VSS.n2667 18.4216
R1258 VSS.n2674 VSS.n2669 18.4216
R1259 VSS.n2670 VSS.n2669 18.4216
R1260 VSS.n2882 VSS.n263 18.4216
R1261 VSS.n2886 VSS.n263 18.4216
R1262 VSS.n2886 VSS.n261 18.4216
R1263 VSS.n2890 VSS.n261 18.4216
R1264 VSS.n2890 VSS.n259 18.4216
R1265 VSS.n2894 VSS.n259 18.4216
R1266 VSS.n2894 VSS.n257 18.4216
R1267 VSS.n2898 VSS.n257 18.4216
R1268 VSS.n2898 VSS.n254 18.4216
R1269 VSS.n2903 VSS.n254 18.4216
R1270 VSS.n2903 VSS.n252 18.4216
R1271 VSS.n2907 VSS.n252 18.4216
R1272 VSS.n2907 VSS.n250 18.4216
R1273 VSS.n2911 VSS.n250 18.4216
R1274 VSS.n2911 VSS.n248 18.4216
R1275 VSS.n2915 VSS.n248 18.4216
R1276 VSS.n2915 VSS.n245 18.4216
R1277 VSS.n2942 VSS.n245 18.4216
R1278 VSS.n2938 VSS.n2927 18.4216
R1279 VSS.n2934 VSS.n2927 18.4216
R1280 VSS.n2934 VSS.n2929 18.4216
R1281 VSS.n2930 VSS.n2929 18.4216
R1282 VSS.n2930 VSS.n200 18.4216
R1283 VSS.n2964 VSS.n200 18.4216
R1284 VSS.n2964 VSS.n198 18.4216
R1285 VSS.n2969 VSS.n198 18.4216
R1286 VSS.n2969 VSS.n196 18.4216
R1287 VSS.n2973 VSS.n196 18.4216
R1288 VSS.n2973 VSS.n193 18.4216
R1289 VSS.n2977 VSS.n193 18.4216
R1290 VSS.n2977 VSS.n191 18.4216
R1291 VSS.n2981 VSS.n191 18.4216
R1292 VSS.n2981 VSS.n189 18.4216
R1293 VSS.n2985 VSS.n189 18.4216
R1294 VSS.n2985 VSS.n187 18.4216
R1295 VSS.n2989 VSS.n187 18.4216
R1296 VSS.n3039 VSS.n173 18.4216
R1297 VSS.n3035 VSS.n173 18.4216
R1298 VSS.n3035 VSS.n2993 18.4216
R1299 VSS.n3031 VSS.n2993 18.4216
R1300 VSS.n3031 VSS.n2994 18.4216
R1301 VSS.n3027 VSS.n2994 18.4216
R1302 VSS.n3027 VSS.n2996 18.4216
R1303 VSS.n3023 VSS.n2996 18.4216
R1304 VSS.n3023 VSS.n2999 18.4216
R1305 VSS.n3019 VSS.n2999 18.4216
R1306 VSS.n3019 VSS.n3001 18.4216
R1307 VSS.n3015 VSS.n3001 18.4216
R1308 VSS.n3015 VSS.n3003 18.4216
R1309 VSS.n3011 VSS.n3003 18.4216
R1310 VSS.n3011 VSS.n3005 18.4216
R1311 VSS.n3007 VSS.n3005 18.4216
R1312 VSS.n3007 VSS.n3 18.4216
R1313 VSS.n3482 VSS.n3 18.4216
R1314 VSS.n327 VSS.n321 18.4216
R1315 VSS.n352 VSS.n318 18.4216
R1316 VSS.n352 VSS.n319 18.4216
R1317 VSS.n348 VSS.n347 18.4216
R1318 VSS.n344 VSS.n343 18.4216
R1319 VSS.n340 VSS.n339 18.4216
R1320 VSS.n336 VSS.n335 18.4216
R1321 VSS.n332 VSS.n331 18.4216
R1322 VSS.n1948 VSS.n1947 18.4216
R1323 VSS.n1945 VSS.n1914 18.4216
R1324 VSS.n1941 VSS.n1914 18.4216
R1325 VSS.n1939 VSS.n1938 18.4216
R1326 VSS.n1936 VSS.n1917 18.4216
R1327 VSS.n1932 VSS.n1931 18.4216
R1328 VSS.n1929 VSS.n1920 18.4216
R1329 VSS.n1925 VSS.n1924 18.4216
R1330 VSS.n1888 VSS.n1887 18.4216
R1331 VSS.n1885 VSS.n1853 18.4216
R1332 VSS.n1881 VSS.n1853 18.4216
R1333 VSS.n1879 VSS.n1878 18.4216
R1334 VSS.n1876 VSS.n1856 18.4216
R1335 VSS.n1872 VSS.n1871 18.4216
R1336 VSS.n1869 VSS.n1859 18.4216
R1337 VSS.n1865 VSS.n1864 18.4216
R1338 VSS.n1809 VSS.n1807 18.4216
R1339 VSS.n1805 VSS.n1773 18.4216
R1340 VSS.n1801 VSS.n1773 18.4216
R1341 VSS.n1799 VSS.n1798 18.4216
R1342 VSS.n1796 VSS.n1776 18.4216
R1343 VSS.n1792 VSS.n1791 18.4216
R1344 VSS.n1789 VSS.n1779 18.4216
R1345 VSS.n1785 VSS.n1784 18.4216
R1346 VSS.n2058 VSS.n2054 18.4216
R1347 VSS.n2089 VSS.n2055 18.4216
R1348 VSS.n2085 VSS.n2055 18.4216
R1349 VSS.n2083 VSS.n2082 18.4216
R1350 VSS.n2080 VSS.n2063 18.4216
R1351 VSS.n2076 VSS.n2075 18.4216
R1352 VSS.n2073 VSS.n2066 18.4216
R1353 VSS.n2069 VSS.n2068 18.4216
R1354 VSS.n2129 VSS.n1771 18.4216
R1355 VSS.n2125 VSS.n1771 18.4216
R1356 VSS.n2125 VSS.n1814 18.4216
R1357 VSS.n2121 VSS.n1814 18.4216
R1358 VSS.n2121 VSS.n1817 18.4216
R1359 VSS.n2117 VSS.n1817 18.4216
R1360 VSS.n2117 VSS.n1819 18.4216
R1361 VSS.n2113 VSS.n1819 18.4216
R1362 VSS.n2113 VSS.n1821 18.4216
R1363 VSS.n2109 VSS.n1821 18.4216
R1364 VSS.n2109 VSS.n1823 18.4216
R1365 VSS.n2105 VSS.n1823 18.4216
R1366 VSS.n2105 VSS.n1825 18.4216
R1367 VSS.n2101 VSS.n1825 18.4216
R1368 VSS.n2101 VSS.n1827 18.4216
R1369 VSS.n2097 VSS.n1827 18.4216
R1370 VSS.n2097 VSS.n1829 18.4216
R1371 VSS.n2093 VSS.n1829 18.4216
R1372 VSS.n2051 VSS.n1831 18.4216
R1373 VSS.n2047 VSS.n1831 18.4216
R1374 VSS.n2047 VSS.n1834 18.4216
R1375 VSS.n2043 VSS.n1834 18.4216
R1376 VSS.n2043 VSS.n1837 18.4216
R1377 VSS.n2039 VSS.n1837 18.4216
R1378 VSS.n2039 VSS.n1839 18.4216
R1379 VSS.n2035 VSS.n1839 18.4216
R1380 VSS.n2035 VSS.n1841 18.4216
R1381 VSS.n2031 VSS.n1841 18.4216
R1382 VSS.n2031 VSS.n1843 18.4216
R1383 VSS.n2027 VSS.n1843 18.4216
R1384 VSS.n2027 VSS.n1845 18.4216
R1385 VSS.n2023 VSS.n1845 18.4216
R1386 VSS.n2023 VSS.n1847 18.4216
R1387 VSS.n2019 VSS.n1847 18.4216
R1388 VSS.n2019 VSS.n1849 18.4216
R1389 VSS.n2015 VSS.n1849 18.4216
R1390 VSS.n2011 VSS.n2010 18.4216
R1391 VSS.n2010 VSS.n1893 18.4216
R1392 VSS.n2006 VSS.n1893 18.4216
R1393 VSS.n2006 VSS.n1895 18.4216
R1394 VSS.n2002 VSS.n1895 18.4216
R1395 VSS.n2002 VSS.n1898 18.4216
R1396 VSS.n1998 VSS.n1898 18.4216
R1397 VSS.n1998 VSS.n1900 18.4216
R1398 VSS.n1994 VSS.n1900 18.4216
R1399 VSS.n1994 VSS.n1902 18.4216
R1400 VSS.n1990 VSS.n1902 18.4216
R1401 VSS.n1990 VSS.n1904 18.4216
R1402 VSS.n1986 VSS.n1904 18.4216
R1403 VSS.n1986 VSS.n1906 18.4216
R1404 VSS.n1982 VSS.n1906 18.4216
R1405 VSS.n1982 VSS.n1908 18.4216
R1406 VSS.n1978 VSS.n1908 18.4216
R1407 VSS.n1978 VSS.n1975 18.4216
R1408 VSS.n1973 VSS.n1911 18.4216
R1409 VSS.n1969 VSS.n1911 18.4216
R1410 VSS.n1969 VSS.n1953 18.4216
R1411 VSS.n1965 VSS.n1953 18.4216
R1412 VSS.n1965 VSS.n1956 18.4216
R1413 VSS.n1961 VSS.n1956 18.4216
R1414 VSS.n1961 VSS.n1958 18.4216
R1415 VSS.n1958 VSS.n83 18.4216
R1416 VSS.n3156 VSS.n83 18.4216
R1417 VSS.n3156 VSS.n84 18.4216
R1418 VSS.n3152 VSS.n84 18.4216
R1419 VSS.n3152 VSS.n87 18.4216
R1420 VSS.n3148 VSS.n87 18.4216
R1421 VSS.n3148 VSS.n90 18.4216
R1422 VSS.n3144 VSS.n90 18.4216
R1423 VSS.n3144 VSS.n92 18.4216
R1424 VSS.n3140 VSS.n92 18.4216
R1425 VSS.n3140 VSS.n94 18.4216
R1426 VSS.n3135 VSS.n98 18.4216
R1427 VSS.n3131 VSS.n98 18.4216
R1428 VSS.n3131 VSS.n101 18.4216
R1429 VSS.n3127 VSS.n101 18.4216
R1430 VSS.n3127 VSS.n103 18.4216
R1431 VSS.n3123 VSS.n103 18.4216
R1432 VSS.n3123 VSS.n105 18.4216
R1433 VSS.n3119 VSS.n105 18.4216
R1434 VSS.n3119 VSS.n107 18.4216
R1435 VSS.n3115 VSS.n107 18.4216
R1436 VSS.n3115 VSS.n108 18.4216
R1437 VSS.n3111 VSS.n108 18.4216
R1438 VSS.n3111 VSS.n110 18.4216
R1439 VSS.n3107 VSS.n110 18.4216
R1440 VSS.n3107 VSS.n113 18.4216
R1441 VSS.n3103 VSS.n113 18.4216
R1442 VSS.n3103 VSS.n115 18.4216
R1443 VSS.n744 VSS.n115 18.4216
R1444 VSS.n748 VSS.n699 18.4216
R1445 VSS.n752 VSS.n699 18.4216
R1446 VSS.n752 VSS.n697 18.4216
R1447 VSS.n756 VSS.n697 18.4216
R1448 VSS.n759 VSS.n758 18.4216
R1449 VSS.n761 VSS.n759 18.4216
R1450 VSS.n765 VSS.n694 18.4216
R1451 VSS.n766 VSS.n765 18.4216
R1452 VSS.n768 VSS.n692 18.4216
R1453 VSS.n772 VSS.n692 18.4216
R1454 VSS.n776 VSS.n774 18.4216
R1455 VSS.n780 VSS.n690 18.4216
R1456 VSS.n913 VSS.n687 18.4216
R1457 VSS.n917 VSS.n915 18.4216
R1458 VSS.n921 VSS.n685 18.4216
R1459 VSS.n925 VSS.n923 18.4216
R1460 VSS.n929 VSS.n683 18.4216
R1461 VSS.n933 VSS.n931 18.4216
R1462 VSS.n937 VSS.n681 18.4216
R1463 VSS.n941 VSS.n939 18.4216
R1464 VSS.n945 VSS.n679 18.4216
R1465 VSS.n739 VSS.n738 18.4216
R1466 VSS.n736 VSS.n704 18.4216
R1467 VSS.n732 VSS.n704 18.4216
R1468 VSS.n730 VSS.n729 18.4216
R1469 VSS.n727 VSS.n707 18.4216
R1470 VSS.n723 VSS.n722 18.4216
R1471 VSS.n720 VSS.n710 18.4216
R1472 VSS.n716 VSS.n715 18.4216
R1473 VSS.n219 VSS.n216 18.4216
R1474 VSS.n222 VSS.n221 18.4216
R1475 VSS.n225 VSS.n222 18.4216
R1476 VSS.n225 VSS.n211 18.4216
R1477 VSS.n229 VSS.n211 18.4216
R1478 VSS.n229 VSS.n209 18.4216
R1479 VSS.n233 VSS.n209 18.4216
R1480 VSS.n233 VSS.n206 18.4216
R1481 VSS.n2958 VSS.n206 18.4216
R1482 VSS.n2958 VSS.n207 18.4216
R1483 VSS.n2954 VSS.n207 18.4216
R1484 VSS.n2954 VSS.n237 18.4216
R1485 VSS.n2950 VSS.n237 18.4216
R1486 VSS.n2950 VSS.n239 18.4216
R1487 VSS.n2946 VSS.n239 18.4216
R1488 VSS.n2946 VSS.n241 18.4216
R1489 VSS.n2922 VSS.n2921 18.4216
R1490 VSS.n2212 VSS.n586 18.4216
R1491 VSS.n2218 VSS.n586 18.4216
R1492 VSS.n2218 VSS.n584 18.4216
R1493 VSS.n2222 VSS.n584 18.4216
R1494 VSS.n2222 VSS.n582 18.4216
R1495 VSS.n2226 VSS.n582 18.4216
R1496 VSS.n2226 VSS.n580 18.4216
R1497 VSS.n2230 VSS.n580 18.4216
R1498 VSS.n2230 VSS.n578 18.4216
R1499 VSS.n2234 VSS.n578 18.4216
R1500 VSS.n2234 VSS.n576 18.4216
R1501 VSS.n2238 VSS.n576 18.4216
R1502 VSS.n2238 VSS.n574 18.4216
R1503 VSS.n2242 VSS.n574 18.4216
R1504 VSS.n2242 VSS.n572 18.4216
R1505 VSS.n2246 VSS.n572 18.4216
R1506 VSS.n2246 VSS.n570 18.4216
R1507 VSS.n2250 VSS.n570 18.4216
R1508 VSS.n2300 VSS.n559 18.4216
R1509 VSS.n2296 VSS.n559 18.4216
R1510 VSS.n2296 VSS.n2254 18.4216
R1511 VSS.n2292 VSS.n2254 18.4216
R1512 VSS.n2292 VSS.n2256 18.4216
R1513 VSS.n2288 VSS.n2256 18.4216
R1514 VSS.n2288 VSS.n2258 18.4216
R1515 VSS.n2284 VSS.n2258 18.4216
R1516 VSS.n2284 VSS.n2260 18.4216
R1517 VSS.n2280 VSS.n2260 18.4216
R1518 VSS.n2280 VSS.n2262 18.4216
R1519 VSS.n2276 VSS.n2262 18.4216
R1520 VSS.n2276 VSS.n2264 18.4216
R1521 VSS.n2272 VSS.n2264 18.4216
R1522 VSS.n2272 VSS.n2266 18.4216
R1523 VSS.n2268 VSS.n2266 18.4216
R1524 VSS.n2268 VSS.n471 18.4216
R1525 VSS.n2472 VSS.n471 18.4216
R1526 VSS.n2476 VSS.n465 18.4216
R1527 VSS.n2480 VSS.n465 18.4216
R1528 VSS.n2480 VSS.n463 18.4216
R1529 VSS.n2484 VSS.n463 18.4216
R1530 VSS.n2484 VSS.n461 18.4216
R1531 VSS.n2488 VSS.n461 18.4216
R1532 VSS.n2488 VSS.n459 18.4216
R1533 VSS.n2492 VSS.n459 18.4216
R1534 VSS.n2492 VSS.n457 18.4216
R1535 VSS.n2496 VSS.n457 18.4216
R1536 VSS.n2496 VSS.n455 18.4216
R1537 VSS.n2500 VSS.n455 18.4216
R1538 VSS.n2500 VSS.n453 18.4216
R1539 VSS.n2504 VSS.n453 18.4216
R1540 VSS.n2504 VSS.n451 18.4216
R1541 VSS.n2508 VSS.n451 18.4216
R1542 VSS.n2508 VSS.n449 18.4216
R1543 VSS.n2512 VSS.n449 18.4216
R1544 VSS.n2567 VSS.n438 18.4216
R1545 VSS.n2563 VSS.n438 18.4216
R1546 VSS.n2563 VSS.n2516 18.4216
R1547 VSS.n2559 VSS.n2516 18.4216
R1548 VSS.n2559 VSS.n2518 18.4216
R1549 VSS.n2555 VSS.n2518 18.4216
R1550 VSS.n2555 VSS.n2520 18.4216
R1551 VSS.n2551 VSS.n2520 18.4216
R1552 VSS.n2551 VSS.n2522 18.4216
R1553 VSS.n2547 VSS.n2522 18.4216
R1554 VSS.n2547 VSS.n2524 18.4216
R1555 VSS.n2543 VSS.n2524 18.4216
R1556 VSS.n2543 VSS.n2526 18.4216
R1557 VSS.n2539 VSS.n2526 18.4216
R1558 VSS.n2539 VSS.n2528 18.4216
R1559 VSS.n2535 VSS.n2528 18.4216
R1560 VSS.n2535 VSS.n2530 18.4216
R1561 VSS.n2531 VSS.n2530 18.4216
R1562 VSS.n2750 VSS.n310 18.4216
R1563 VSS.n2750 VSS.n308 18.4216
R1564 VSS.n2754 VSS.n308 18.4216
R1565 VSS.n2754 VSS.n306 18.4216
R1566 VSS.n2758 VSS.n306 18.4216
R1567 VSS.n2758 VSS.n304 18.4216
R1568 VSS.n2762 VSS.n304 18.4216
R1569 VSS.n2762 VSS.n302 18.4216
R1570 VSS.n2766 VSS.n302 18.4216
R1571 VSS.n2766 VSS.n300 18.4216
R1572 VSS.n2770 VSS.n300 18.4216
R1573 VSS.n2770 VSS.n298 18.4216
R1574 VSS.n2774 VSS.n298 18.4216
R1575 VSS.n2774 VSS.n296 18.4216
R1576 VSS.n2779 VSS.n296 18.4216
R1577 VSS.n2779 VSS.n294 18.4216
R1578 VSS.n2783 VSS.n294 18.4216
R1579 VSS.n2784 VSS.n2783 18.4216
R1580 VSS.n2832 VSS.n2787 18.4216
R1581 VSS.n2828 VSS.n2787 18.4216
R1582 VSS.n2828 VSS.n2789 18.4216
R1583 VSS.n2824 VSS.n2789 18.4216
R1584 VSS.n2824 VSS.n2791 18.4216
R1585 VSS.n2820 VSS.n2791 18.4216
R1586 VSS.n2820 VSS.n2793 18.4216
R1587 VSS.n2816 VSS.n2793 18.4216
R1588 VSS.n2816 VSS.n2795 18.4216
R1589 VSS.n2812 VSS.n2795 18.4216
R1590 VSS.n2812 VSS.n2797 18.4216
R1591 VSS.n2808 VSS.n2797 18.4216
R1592 VSS.n2808 VSS.n2799 18.4216
R1593 VSS.n2804 VSS.n2799 18.4216
R1594 VSS.n2804 VSS.n2801 18.4216
R1595 VSS.n2801 VSS.n120 18.4216
R1596 VSS.n3099 VSS.n120 18.4216
R1597 VSS.n3099 VSS.n121 18.4216
R1598 VSS.n3094 VSS.n127 18.4216
R1599 VSS.n3090 VSS.n127 18.4216
R1600 VSS.n3090 VSS.n131 18.4216
R1601 VSS.n3086 VSS.n131 18.4216
R1602 VSS.n3084 VSS.n3083 18.4216
R1603 VSS.n3081 VSS.n135 18.4216
R1604 VSS.n3077 VSS.n135 18.4216
R1605 VSS.n3077 VSS.n137 18.4216
R1606 VSS.n3073 VSS.n137 18.4216
R1607 VSS.n3073 VSS.n144 18.4216
R1608 VSS.n3069 VSS.n144 18.4216
R1609 VSS.n3069 VSS.n146 18.4216
R1610 VSS.n3065 VSS.n146 18.4216
R1611 VSS.n3065 VSS.n148 18.4216
R1612 VSS.n3061 VSS.n148 18.4216
R1613 VSS.n3061 VSS.n150 18.4216
R1614 VSS.n886 VSS.n796 18.4216
R1615 VSS.n882 VSS.n796 18.4216
R1616 VSS.n882 VSS.n834 18.4216
R1617 VSS.n878 VSS.n834 18.4216
R1618 VSS.n878 VSS.n835 18.4216
R1619 VSS.n874 VSS.n835 18.4216
R1620 VSS.n874 VSS.n837 18.4216
R1621 VSS.n870 VSS.n837 18.4216
R1622 VSS.n870 VSS.n840 18.4216
R1623 VSS.n866 VSS.n840 18.4216
R1624 VSS.n866 VSS.n863 18.4216
R1625 VSS.n863 VSS.n862 18.4216
R1626 VSS.n862 VSS.n842 18.4216
R1627 VSS.n858 VSS.n857 18.4216
R1628 VSS.n855 VSS.n845 18.4216
R1629 VSS.n906 VSS.n783 18.4216
R1630 VSS.n902 VSS.n783 18.4216
R1631 VSS.n902 VSS.n786 18.4216
R1632 VSS.n898 VSS.n786 18.4216
R1633 VSS.n898 VSS.n896 18.4216
R1634 VSS.n894 VSS.n790 18.4216
R1635 VSS.n890 VSS.n790 18.4216
R1636 VSS.n890 VSS.n792 18.4216
R1637 VSS.n801 VSS.n792 18.4216
R1638 VSS.n805 VSS.n803 18.4216
R1639 VSS.n809 VSS.n798 18.4216
R1640 VSS.n812 VSS.n811 18.4216
R1641 VSS.n2303 VSS.n552 17.4841
R1642 VSS.n2470 VSS.n476 17.4841
R1643 VSS.n2570 VSS.n432 17.4841
R1644 VSS.n2746 VSS.n2745 17.4841
R1645 VSS.n2842 VSS.n2841 17.4841
R1646 VSS.n1346 VSS.n1226 16.9479
R1647 VSS.n1310 VSS.n1227 16.9479
R1648 VSS.n1360 VSS.n1351 16.5247
R1649 VSS.n322 VSS.n93 16.1749
R1650 VSS.n111 VSS.t17 16.1749
R1651 VSS.t320 VSS.t96 15.6666
R1652 VSS.n1640 VSS.n1083 14.5036
R1653 VSS.n849 VSS.n38 14.142
R1654 VSS.n1252 VSS.n1251 13.8958
R1655 VSS.n3446 VSS.n39 13.706
R1656 VSS.n1650 VSS.n1649 13.676
R1657 VSS.n1627 VSS.n1626 13.5743
R1658 VSS.n949 VSS.n948 13.0685
R1659 VSS.t18 VSS.n1959 12.9931
R1660 VSS.n2300 VSS.n558 12.5268
R1661 VSS.n2476 VSS.n467 12.5268
R1662 VSS.n2567 VSS.n437 12.5268
R1663 VSS.n360 VSS.n310 12.5268
R1664 VSS.n2832 VSS.n290 12.5268
R1665 VSS.n3094 VSS.n126 12.5268
R1666 VSS.n886 VSS.n795 12.5268
R1667 VSS.n2155 VSS.n613 12.4628
R1668 VSS.n325 VSS.n322 12.4628
R1669 VSS.n1513 VSS.t213 12.4059
R1670 VSS.n2360 VSS.t261 12.4059
R1671 VSS.n2394 VSS.t228 12.4059
R1672 VSS.n2627 VSS.t265 12.4059
R1673 VSS.n2661 VSS.t263 12.4059
R1674 VSS.n255 VSS.t211 12.4059
R1675 VSS.n194 VSS.t283 12.3005
R1676 VSS.n1581 VSS.n1575 12.033
R1677 VSS.n1581 VSS.n1574 12.033
R1678 VSS.n1431 VSS.n1418 12.033
R1679 VSS.n3444 VSS.t313 11.9233
R1680 VSS.n2997 VSS.n159 11.6366
R1681 VSS.n21 VSS.n15 11.4244
R1682 VSS.n2345 VSS.n529 11.4216
R1683 VSS.n2435 VSS.n498 11.4216
R1684 VSS.n2612 VSS.n409 11.4216
R1685 VSS.n2707 VSS.n380 11.4216
R1686 VSS.n2882 VSS.n265 11.4216
R1687 VSS.n2938 VSS.n246 11.4216
R1688 VSS.n3039 VSS.n172 11.4216
R1689 VSS.n2052 VSS.n2051 11.4216
R1690 VSS.n2011 VSS.n1850 11.4216
R1691 VSS.n1974 VSS.n1973 11.4216
R1692 VSS.n3135 VSS.n97 11.4216
R1693 VSS.n748 VSS.n701 11.4216
R1694 VSS.n909 VSS.n907 11.4216
R1695 VSS.n3479 VSS.n3478 11.3366
R1696 VSS.n677 VSS.t160 11.1395
R1697 VSS.n1580 VSS.t298 11.0292
R1698 VSS.n1580 VSS.t152 11.0292
R1699 VSS.n1433 VSS.t119 11.0292
R1700 VSS.n1151 VSS.t155 11.0225
R1701 VSS.n3450 VSS.n38 10.6136
R1702 VSS.t183 VSS.n3157 10.6067
R1703 VSS.n1598 VSS.t230 10.5091
R1704 VSS.n3429 VSS.n3159 10.4005
R1705 VSS.n3429 VSS.n78 10.4005
R1706 VSS.n3429 VSS.n3160 10.4005
R1707 VSS.n3429 VSS.n77 10.4005
R1708 VSS.n3429 VSS.n3161 10.4005
R1709 VSS.n3429 VSS.n76 10.4005
R1710 VSS.n3429 VSS.n3162 10.4005
R1711 VSS.n3429 VSS.n75 10.4005
R1712 VSS.n3429 VSS.n3163 10.4005
R1713 VSS.n3429 VSS.n74 10.4005
R1714 VSS.n3429 VSS.n3164 10.4005
R1715 VSS.n3429 VSS.n73 10.4005
R1716 VSS.n3429 VSS.n3165 10.4005
R1717 VSS.n3429 VSS.n72 10.4005
R1718 VSS.n3429 VSS.n3428 10.4005
R1719 VSS.n3429 VSS.n71 10.4005
R1720 VSS.n3430 VSS.n3429 10.4005
R1721 VSS.n1388 VSS.n1387 10.4005
R1722 VSS.n1385 VSS.n1384 10.4005
R1723 VSS.n1153 VSS.n1152 10.4005
R1724 VSS.n1381 VSS.n1380 10.4005
R1725 VSS.n1154 VSS.t154 10.4005
R1726 VSS.t42 VSS.n1383 10.4005
R1727 VSS.n1382 VSS.t71 10.4005
R1728 VSS.t68 VSS.n1155 10.4005
R1729 VSS.n1651 VSS.n1650 10.4005
R1730 VSS.n1626 VSS.n1625 10.4005
R1731 VSS.n1621 VSS.n1094 10.3255
R1732 VSS.n1408 VSS.t240 10.2792
R1733 VSS.n1566 VSS.t242 10.2607
R1734 VSS.n1597 VSS.t53 10.0514
R1735 VSS.n1595 VSS.t57 10.0514
R1736 VSS.t291 VSS.t63 9.96983
R1737 VSS.n1245 VSS.n1244 9.94787
R1738 VSS.n1250 VSS.n1249 9.94787
R1739 VSS.n2341 VSS.n529 9.94787
R1740 VSS.n2383 VSS.n498 9.94787
R1741 VSS.n2608 VSS.n409 9.94787
R1742 VSS.n2650 VSS.n380 9.94787
R1743 VSS.n2670 VSS.n265 9.94787
R1744 VSS.n2942 VSS.n246 9.94787
R1745 VSS.n2989 VSS.n172 9.94787
R1746 VSS.n2093 VSS.n2052 9.94787
R1747 VSS.n2015 VSS.n1850 9.94787
R1748 VSS.n1975 VSS.n1974 9.94787
R1749 VSS.n97 VSS.n94 9.94787
R1750 VSS.n744 VSS.n701 9.94787
R1751 VSS.n907 VSS.n782 9.94787
R1752 VSS.n1144 VSS.t73 9.93604
R1753 VSS.n1140 VSS.t24 9.93604
R1754 VSS.n1137 VSS.t35 9.93604
R1755 VSS.n1127 VSS.t178 9.93604
R1756 VSS.n1422 VSS.t182 9.93604
R1757 VSS.n1428 VSS.t65 9.93604
R1758 VSS.n1429 VSS.t305 9.93604
R1759 VSS.n1437 VSS.t301 9.93604
R1760 VSS.n1437 VSS.t300 9.93604
R1761 VSS.t280 VSS.t165 9.87463
R1762 VSS.n1619 VSS.t28 9.84591
R1763 VSS.n1554 VSS.n1407 9.73801
R1764 VSS.n2303 VSS.n2302 9.71359
R1765 VSS.n476 VSS.n466 9.71359
R1766 VSS.n2570 VSS.n2569 9.71359
R1767 VSS.n2747 VSS.n2746 9.71359
R1768 VSS.n2842 VSS.n99 9.71359
R1769 VSS.n849 VSS.n25 9.19675
R1770 VSS.n3465 VSS.n21 9.188
R1771 VSS.n1594 VSS.t312 9.15882
R1772 VSS.n29 VSS.t333 9.05408
R1773 VSS.n2212 VSS.n592 9.02682
R1774 VSS.n1381 VSS.t68 9.01367
R1775 VSS.n3444 VSS.n3443 8.92063
R1776 VSS.n2250 VSS.n558 8.84261
R1777 VSS.n2472 VSS.n467 8.84261
R1778 VSS.n2512 VSS.n437 8.84261
R1779 VSS.n2531 VSS.n360 8.84261
R1780 VSS.n2784 VSS.n290 8.84261
R1781 VSS.n126 VSS.n121 8.84261
R1782 VSS.n795 VSS.n150 8.84261
R1783 VSS.n3432 VSS.n68 8.77991
R1784 VSS.n1395 VSS.t126 8.51132
R1785 VSS.n1396 VSS.t61 8.51132
R1786 VSS.n1399 VSS.t279 8.51132
R1787 VSS.n1616 VSS.t176 8.51132
R1788 VSS.n1570 VSS.t30 8.51132
R1789 VSS.n1578 VSS.t44 8.51132
R1790 VSS.n1578 VSS.t76 8.51132
R1791 VSS.n1081 VSS.t105 8.51132
R1792 VSS.n1084 VSS.t218 8.51132
R1793 VSS.n1085 VSS.t48 8.51132
R1794 VSS.n1086 VSS.t252 8.51132
R1795 VSS.n1087 VSS.t97 8.51132
R1796 VSS.n1111 VSS.t180 8.51132
R1797 VSS.n1112 VSS.t185 8.51132
R1798 VSS.n1114 VSS.t348 8.51132
R1799 VSS.n1115 VSS.t95 8.51132
R1800 VSS.n1128 VSS.t163 8.51132
R1801 VSS.n1130 VSS.t91 8.51132
R1802 VSS.n1132 VSS.t215 8.51132
R1803 VSS.n1133 VSS.t297 8.51132
R1804 VSS.n1135 VSS.t128 8.51132
R1805 VSS.n1138 VSS.t22 8.51132
R1806 VSS.n1421 VSS.t16 8.51132
R1807 VSS.n1569 VSS.t111 8.51132
R1808 VSS.n1141 VSS.t303 8.48197
R1809 VSS.n1583 VSS.t11 8.46241
R1810 VSS.n1583 VSS.t130 8.46241
R1811 VSS.n1425 VSS.t342 8.46241
R1812 VSS.n1142 VSS.t78 8.4135
R1813 VSS.n1134 VSS.t327 8.4135
R1814 VSS.n1131 VSS.t32 8.4135
R1815 VSS.n1129 VSS.t310 8.4135
R1816 VSS.n1426 VSS.t132 8.4135
R1817 VSS.n1432 VSS.t234 8.4135
R1818 VSS.n1434 VSS.t307 8.4135
R1819 VSS.n1436 VSS.t70 8.4135
R1820 VSS.n1575 VSS.t79 8.4005
R1821 VSS.n1575 VSS.t41 8.4005
R1822 VSS.n1574 VSS.t13 8.4005
R1823 VSS.n1574 VSS.t85 8.4005
R1824 VSS.n1418 VSS.t39 8.4005
R1825 VSS.n1418 VSS.t124 8.4005
R1826 VSS.n2130 VSS.n2129 8.14755
R1827 VSS.n1573 VSS.t9 8.0855
R1828 VSS.n1572 VSS.t129 8.0855
R1829 VSS.n1420 VSS.t340 8.0855
R1830 VSS.n534 VSS.n529 7.92155
R1831 VSS.n508 VSS.n498 7.92155
R1832 VSS.n414 VSS.n409 7.92155
R1833 VSS.n388 VSS.n380 7.92155
R1834 VSS.n2871 VSS.n265 7.92155
R1835 VSS.n184 VSS.n172 7.92155
R1836 VSS.n2924 VSS.n246 7.92155
R1837 VSS.n566 VSS.n558 7.82945
R1838 VSS.n477 VSS.n467 7.82945
R1839 VSS.n445 VSS.n437 7.82945
R1840 VSS.n2743 VSS.n360 7.82945
R1841 VSS.n2839 VSS.n290 7.82945
R1842 VSS.n830 VSS.n795 7.82945
R1843 VSS.n214 VSS.n126 7.82945
R1844 VSS.n1247 VSS.n1218 7.74316
R1845 VSS.n1262 VSS.n1226 7.36892
R1846 VSS.n1310 VSS.n1309 7.36892
R1847 VSS.n1241 VSS.t2 7.13593
R1848 VSS.n1248 VSS.t0 7.13593
R1849 VSS.n1097 VSS.t147 7.06906
R1850 VSS.n1352 VSS.n1091 6.94217
R1851 VSS.n3101 VSS.n116 6.62937
R1852 VSS.n15 VSS.n4 6.62351
R1853 VSS.n1582 VSS.n1572 6.54898
R1854 VSS.n1582 VSS.n1573 6.54898
R1855 VSS.n1427 VSS.n1420 6.54898
R1856 VSS.n1398 VSS.n1397 6.50202
R1857 VSS.n1101 VSS.n1100 6.50202
R1858 VSS.n1615 VSS.n1099 6.50202
R1859 VSS.n1618 VSS.n1097 6.4805
R1860 VSS.n1579 VSS.n1576 6.46859
R1861 VSS.n1579 VSS.n1577 6.46859
R1862 VSS.n1435 VSS.n1417 6.46859
R1863 VSS.n1599 VSS.n1409 6.46462
R1864 VSS.n1565 VSS.n1560 6.45138
R1865 VSS.n1564 VSS.n1561 6.45138
R1866 VSS.n1563 VSS.n1562 6.45138
R1867 VSS.n1596 VSS.n1410 6.45138
R1868 VSS.n323 VSS.n97 6.44787
R1869 VSS.n1974 VSS.n1910 6.44787
R1870 VSS.n1890 VSS.n1850 6.44787
R1871 VSS.n2130 VSS.n1770 6.44787
R1872 VSS.n2056 VSS.n2052 6.44787
R1873 VSS.n946 VSS.n945 6.44787
R1874 VSS.n741 VSS.n701 6.44787
R1875 VSS.n907 VSS.n906 6.44787
R1876 VSS.n1110 VSS.t62 6.3005
R1877 VSS.n851 VSS.n850 6.17155
R1878 VSS.n1388 VSS.t154 6.00928
R1879 VSS.n2215 VSS.n2214 5.82835
R1880 VSS.n848 VSS.n25 5.63714
R1881 VSS.n1110 VSS.t352 5.6196
R1882 VSS.n2215 VSS.n590 5.5943
R1883 VSS.n678 VSS.n42 5.39487
R1884 VSS.n1644 VSS.n1643 5.32359
R1885 VSS.n1118 VSS.n1117 5.32359
R1886 VSS.n1139 VSS.n1123 5.32359
R1887 VSS.n1143 VSS.n1122 5.32359
R1888 VSS.n1145 VSS.n1121 5.32359
R1889 VSS.n1146 VSS.n1120 5.32359
R1890 VSS.n1424 VSS.n1423 5.32359
R1891 VSS.n1571 VSS.n1559 5.32359
R1892 VSS.n1401 VSS.n1400 5.32226
R1893 VSS.n1585 VSS.n1584 5.32226
R1894 VSS.n1126 VSS.n1125 5.32226
R1895 VSS.n1136 VSS.n1124 5.32226
R1896 VSS.n1430 VSS.n1419 5.32226
R1897 VSS.n1617 VSS.n1098 5.32226
R1898 VSS.n1593 VSS.n1411 5.32226
R1899 VSS.n2997 VSS.n2994 5.23035
R1900 VSS.n1203 VSS.n1163 5.2014
R1901 VSS.n2306 VSS.n2305 5.2005
R1902 VSS.n2305 VSS.n2304 5.2005
R1903 VSS.n2307 VSS.n549 5.2005
R1904 VSS.n549 VSS.n548 5.2005
R1905 VSS.n2309 VSS.n2308 5.2005
R1906 VSS.n2310 VSS.n2309 5.2005
R1907 VSS.n547 VSS.n546 5.2005
R1908 VSS.n2311 VSS.n547 5.2005
R1909 VSS.n2314 VSS.n2313 5.2005
R1910 VSS.n2313 VSS.n2312 5.2005
R1911 VSS.n2315 VSS.n545 5.2005
R1912 VSS.n545 VSS.n544 5.2005
R1913 VSS.n2317 VSS.n2316 5.2005
R1914 VSS.n2318 VSS.n2317 5.2005
R1915 VSS.n543 VSS.n542 5.2005
R1916 VSS.n2319 VSS.n543 5.2005
R1917 VSS.n2322 VSS.n2321 5.2005
R1918 VSS.n2321 VSS.n2320 5.2005
R1919 VSS.n2323 VSS.n541 5.2005
R1920 VSS.n541 VSS.n540 5.2005
R1921 VSS.n2325 VSS.n2324 5.2005
R1922 VSS.n2326 VSS.n2325 5.2005
R1923 VSS.n539 VSS.n538 5.2005
R1924 VSS.n2327 VSS.n539 5.2005
R1925 VSS.n2331 VSS.n2330 5.2005
R1926 VSS.n2330 VSS.n2329 5.2005
R1927 VSS.n2332 VSS.n537 5.2005
R1928 VSS.n2328 VSS.n537 5.2005
R1929 VSS.n2465 VSS.n2464 5.2005
R1930 VSS.n2464 VSS.n2463 5.2005
R1931 VSS.n483 VSS.n482 5.2005
R1932 VSS.n2462 VSS.n483 5.2005
R1933 VSS.n2460 VSS.n2459 5.2005
R1934 VSS.n2461 VSS.n2460 5.2005
R1935 VSS.n2458 VSS.n485 5.2005
R1936 VSS.n485 VSS.n484 5.2005
R1937 VSS.n2457 VSS.n2456 5.2005
R1938 VSS.n2456 VSS.n2455 5.2005
R1939 VSS.n487 VSS.n486 5.2005
R1940 VSS.n2454 VSS.n487 5.2005
R1941 VSS.n2452 VSS.n2451 5.2005
R1942 VSS.n2453 VSS.n2452 5.2005
R1943 VSS.n2450 VSS.n489 5.2005
R1944 VSS.n489 VSS.n488 5.2005
R1945 VSS.n2449 VSS.n2448 5.2005
R1946 VSS.n2448 VSS.n2447 5.2005
R1947 VSS.n491 VSS.n490 5.2005
R1948 VSS.n2446 VSS.n491 5.2005
R1949 VSS.n2444 VSS.n2443 5.2005
R1950 VSS.n2445 VSS.n2444 5.2005
R1951 VSS.n2442 VSS.n493 5.2005
R1952 VSS.n493 VSS.n492 5.2005
R1953 VSS.n2441 VSS.n2440 5.2005
R1954 VSS.n2440 VSS.n2439 5.2005
R1955 VSS.n495 VSS.n494 5.2005
R1956 VSS.n2438 VSS.n495 5.2005
R1957 VSS.n2573 VSS.n2572 5.2005
R1958 VSS.n2572 VSS.n2571 5.2005
R1959 VSS.n2574 VSS.n429 5.2005
R1960 VSS.n429 VSS.n428 5.2005
R1961 VSS.n2576 VSS.n2575 5.2005
R1962 VSS.n2577 VSS.n2576 5.2005
R1963 VSS.n427 VSS.n426 5.2005
R1964 VSS.n2578 VSS.n427 5.2005
R1965 VSS.n2581 VSS.n2580 5.2005
R1966 VSS.n2580 VSS.n2579 5.2005
R1967 VSS.n2582 VSS.n425 5.2005
R1968 VSS.n425 VSS.n424 5.2005
R1969 VSS.n2584 VSS.n2583 5.2005
R1970 VSS.n2585 VSS.n2584 5.2005
R1971 VSS.n423 VSS.n422 5.2005
R1972 VSS.n2586 VSS.n423 5.2005
R1973 VSS.n2589 VSS.n2588 5.2005
R1974 VSS.n2588 VSS.n2587 5.2005
R1975 VSS.n2590 VSS.n421 5.2005
R1976 VSS.n421 VSS.n420 5.2005
R1977 VSS.n2592 VSS.n2591 5.2005
R1978 VSS.n2593 VSS.n2592 5.2005
R1979 VSS.n419 VSS.n418 5.2005
R1980 VSS.n2594 VSS.n419 5.2005
R1981 VSS.n2598 VSS.n2597 5.2005
R1982 VSS.n2597 VSS.n2596 5.2005
R1983 VSS.n2599 VSS.n417 5.2005
R1984 VSS.n2595 VSS.n417 5.2005
R1985 VSS.n2736 VSS.n362 5.2005
R1986 VSS.n2736 VSS.n354 5.2005
R1987 VSS.n2735 VSS.n364 5.2005
R1988 VSS.n2735 VSS.n2734 5.2005
R1989 VSS.n367 VSS.n363 5.2005
R1990 VSS.n2733 VSS.n363 5.2005
R1991 VSS.n2731 VSS.n2730 5.2005
R1992 VSS.n2732 VSS.n2731 5.2005
R1993 VSS.n2729 VSS.n366 5.2005
R1994 VSS.n366 VSS.n365 5.2005
R1995 VSS.n2728 VSS.n2727 5.2005
R1996 VSS.n2727 VSS.n2726 5.2005
R1997 VSS.n369 VSS.n368 5.2005
R1998 VSS.n2725 VSS.n369 5.2005
R1999 VSS.n2723 VSS.n2722 5.2005
R2000 VSS.n2724 VSS.n2723 5.2005
R2001 VSS.n2721 VSS.n371 5.2005
R2002 VSS.n371 VSS.n370 5.2005
R2003 VSS.n2720 VSS.n2719 5.2005
R2004 VSS.n2719 VSS.n2718 5.2005
R2005 VSS.n373 VSS.n372 5.2005
R2006 VSS.n2717 VSS.n373 5.2005
R2007 VSS.n2715 VSS.n2714 5.2005
R2008 VSS.n2716 VSS.n2715 5.2005
R2009 VSS.n2713 VSS.n375 5.2005
R2010 VSS.n375 VSS.n374 5.2005
R2011 VSS.n2712 VSS.n2711 5.2005
R2012 VSS.n2711 VSS.n2710 5.2005
R2013 VSS.n2845 VSS.n2844 5.2005
R2014 VSS.n2844 VSS.n2843 5.2005
R2015 VSS.n2846 VSS.n282 5.2005
R2016 VSS.n282 VSS.n281 5.2005
R2017 VSS.n2848 VSS.n2847 5.2005
R2018 VSS.n2849 VSS.n2848 5.2005
R2019 VSS.n280 VSS.n279 5.2005
R2020 VSS.n2850 VSS.n280 5.2005
R2021 VSS.n2853 VSS.n2852 5.2005
R2022 VSS.n2852 VSS.n2851 5.2005
R2023 VSS.n2854 VSS.n278 5.2005
R2024 VSS.n278 VSS.n277 5.2005
R2025 VSS.n2856 VSS.n2855 5.2005
R2026 VSS.n2857 VSS.n2856 5.2005
R2027 VSS.n276 VSS.n275 5.2005
R2028 VSS.n2858 VSS.n276 5.2005
R2029 VSS.n2861 VSS.n2860 5.2005
R2030 VSS.n2860 VSS.n2859 5.2005
R2031 VSS.n2862 VSS.n274 5.2005
R2032 VSS.n274 VSS.n273 5.2005
R2033 VSS.n2864 VSS.n2863 5.2005
R2034 VSS.n2865 VSS.n2864 5.2005
R2035 VSS.n272 VSS.n271 5.2005
R2036 VSS.n2866 VSS.n272 5.2005
R2037 VSS.n2869 VSS.n2868 5.2005
R2038 VSS.n2868 VSS.n2867 5.2005
R2039 VSS.n2870 VSS.n270 5.2005
R2040 VSS.n270 VSS.n266 5.2005
R2041 VSS.n1885 VSS.n1884 5.2005
R2042 VSS.n1887 VSS.n1852 5.2005
R2043 VSS.n1888 VSS.n1851 5.2005
R2044 VSS.n1891 VSS.n1890 5.2005
R2045 VSS.n1945 VSS.n1944 5.2005
R2046 VSS.n1947 VSS.n1912 5.2005
R2047 VSS.n1949 VSS.n1948 5.2005
R2048 VSS.n1950 VSS.n1910 5.2005
R2049 VSS.n329 VSS.n318 5.2005
R2050 VSS.n328 VSS.n327 5.2005
R2051 VSS.n321 VSS.n320 5.2005
R2052 VSS.n323 VSS.n95 5.2005
R2053 VSS.n1805 VSS.n1804 5.2005
R2054 VSS.n1807 VSS.n1772 5.2005
R2055 VSS.n1810 VSS.n1809 5.2005
R2056 VSS.n1811 VSS.n1770 5.2005
R2057 VSS.n1789 VSS.n1788 5.2005
R2058 VSS.n1791 VSS.n1777 5.2005
R2059 VSS.n1793 VSS.n1792 5.2005
R2060 VSS.n1794 VSS.n1776 5.2005
R2061 VSS.n1796 VSS.n1795 5.2005
R2062 VSS.n1798 VSS.n1775 5.2005
R2063 VSS.n1799 VSS.n1774 5.2005
R2064 VSS.n1802 VSS.n1801 5.2005
R2065 VSS.n1803 VSS.n1773 5.2005
R2066 VSS.n1773 VSS.n555 5.2005
R2067 VSS.n1869 VSS.n1868 5.2005
R2068 VSS.n1871 VSS.n1857 5.2005
R2069 VSS.n1873 VSS.n1872 5.2005
R2070 VSS.n1874 VSS.n1856 5.2005
R2071 VSS.n1876 VSS.n1875 5.2005
R2072 VSS.n1878 VSS.n1855 5.2005
R2073 VSS.n1879 VSS.n1854 5.2005
R2074 VSS.n1882 VSS.n1881 5.2005
R2075 VSS.n1883 VSS.n1853 5.2005
R2076 VSS.n1853 VSS.n435 5.2005
R2077 VSS.n1929 VSS.n1928 5.2005
R2078 VSS.n1931 VSS.n1918 5.2005
R2079 VSS.n1933 VSS.n1932 5.2005
R2080 VSS.n1934 VSS.n1917 5.2005
R2081 VSS.n1936 VSS.n1935 5.2005
R2082 VSS.n1938 VSS.n1916 5.2005
R2083 VSS.n1939 VSS.n1915 5.2005
R2084 VSS.n1942 VSS.n1941 5.2005
R2085 VSS.n1943 VSS.n1914 5.2005
R2086 VSS.n1914 VSS.n313 5.2005
R2087 VSS.n337 VSS.n336 5.2005
R2088 VSS.n339 VSS.n338 5.2005
R2089 VSS.n341 VSS.n340 5.2005
R2090 VSS.n343 VSS.n342 5.2005
R2091 VSS.n345 VSS.n344 5.2005
R2092 VSS.n347 VSS.n346 5.2005
R2093 VSS.n349 VSS.n348 5.2005
R2094 VSS.n350 VSS.n319 5.2005
R2095 VSS.n352 VSS.n351 5.2005
R2096 VSS.n353 VSS.n352 5.2005
R2097 VSS.n3044 VSS.n3043 5.2005
R2098 VSS.n166 VSS.n162 5.2005
R2099 VSS.n175 VSS.n174 5.2005
R2100 VSS.n177 VSS.n176 5.2005
R2101 VSS.n179 VSS.n178 5.2005
R2102 VSS.n181 VSS.n180 5.2005
R2103 VSS.n183 VSS.n182 5.2005
R2104 VSS.n185 VSS.n184 5.2005
R2105 VSS.n2877 VSS.n2876 5.2005
R2106 VSS.n2875 VSS.n269 5.2005
R2107 VSS.n2874 VSS.n2873 5.2005
R2108 VSS.n2872 VSS.n2871 5.2005
R2109 VSS.n377 VSS.n376 5.2005
R2110 VSS.n385 VSS.n383 5.2005
R2111 VSS.n386 VSS.n382 5.2005
R2112 VSS.n389 VSS.n388 5.2005
R2113 VSS.n2604 VSS.n2603 5.2005
R2114 VSS.n2602 VSS.n416 5.2005
R2115 VSS.n2601 VSS.n2600 5.2005
R2116 VSS.n414 VSS.n410 5.2005
R2117 VSS.n503 VSS.n502 5.2005
R2118 VSS.n505 VSS.n501 5.2005
R2119 VSS.n506 VSS.n500 5.2005
R2120 VSS.n509 VSS.n508 5.2005
R2121 VSS.n2337 VSS.n2336 5.2005
R2122 VSS.n2335 VSS.n536 5.2005
R2123 VSS.n2334 VSS.n2333 5.2005
R2124 VSS.n534 VSS.n530 5.2005
R2125 VSS.n2839 VSS.n2838 5.2005
R2126 VSS.n2837 VSS.n289 5.2005
R2127 VSS.n2836 VSS.n2835 5.2005
R2128 VSS.n284 VSS.n283 5.2005
R2129 VSS.n2743 VSS.n2742 5.2005
R2130 VSS.n2741 VSS.n359 5.2005
R2131 VSS.n2740 VSS.n2739 5.2005
R2132 VSS.n2738 VSS.n2737 5.2005
R2133 VSS.n446 VSS.n445 5.2005
R2134 VSS.n443 VSS.n439 5.2005
R2135 VSS.n442 VSS.n441 5.2005
R2136 VSS.n431 VSS.n430 5.2005
R2137 VSS.n477 VSS.n468 5.2005
R2138 VSS.n481 VSS.n480 5.2005
R2139 VSS.n2468 VSS.n2467 5.2005
R2140 VSS.n2466 VSS.n479 5.2005
R2141 VSS.n567 VSS.n566 5.2005
R2142 VSS.n564 VSS.n560 5.2005
R2143 VSS.n563 VSS.n562 5.2005
R2144 VSS.n551 VSS.n550 5.2005
R2145 VSS.n1782 VSS.n568 5.2005
R2146 VSS.n1784 VSS.n1780 5.2005
R2147 VSS.n1786 VSS.n1785 5.2005
R2148 VSS.n1787 VSS.n1779 5.2005
R2149 VSS.n1862 VSS.n447 5.2005
R2150 VSS.n1864 VSS.n1860 5.2005
R2151 VSS.n1866 VSS.n1865 5.2005
R2152 VSS.n1867 VSS.n1859 5.2005
R2153 VSS.n1922 VSS.n1921 5.2005
R2154 VSS.n1924 VSS.n1923 5.2005
R2155 VSS.n1926 VSS.n1925 5.2005
R2156 VSS.n1927 VSS.n1920 5.2005
R2157 VSS.n292 VSS.n291 5.2005
R2158 VSS.n331 VSS.n330 5.2005
R2159 VSS.n333 VSS.n332 5.2005
R2160 VSS.n335 VSS.n334 5.2005
R2161 VSS.n474 VSS.n469 5.2005
R2162 VSS.n2068 VSS.n2067 5.2005
R2163 VSS.n2070 VSS.n2069 5.2005
R2164 VSS.n2071 VSS.n2066 5.2005
R2165 VSS.n2073 VSS.n2072 5.2005
R2166 VSS.n2075 VSS.n2064 5.2005
R2167 VSS.n2077 VSS.n2076 5.2005
R2168 VSS.n2078 VSS.n2063 5.2005
R2169 VSS.n2080 VSS.n2079 5.2005
R2170 VSS.n2082 VSS.n2062 5.2005
R2171 VSS.n2083 VSS.n2061 5.2005
R2172 VSS.n2086 VSS.n2085 5.2005
R2173 VSS.n2087 VSS.n2055 5.2005
R2174 VSS.n2055 VSS.n556 5.2005
R2175 VSS.n2089 VSS.n2088 5.2005
R2176 VSS.n2060 VSS.n2054 5.2005
R2177 VSS.n2059 VSS.n2058 5.2005
R2178 VSS.n2057 VSS.n2056 5.2005
R2179 VSS.n713 VSS.n124 5.2005
R2180 VSS.n715 VSS.n711 5.2005
R2181 VSS.n717 VSS.n716 5.2005
R2182 VSS.n718 VSS.n710 5.2005
R2183 VSS.n720 VSS.n719 5.2005
R2184 VSS.n722 VSS.n708 5.2005
R2185 VSS.n724 VSS.n723 5.2005
R2186 VSS.n725 VSS.n707 5.2005
R2187 VSS.n727 VSS.n726 5.2005
R2188 VSS.n729 VSS.n706 5.2005
R2189 VSS.n730 VSS.n705 5.2005
R2190 VSS.n733 VSS.n732 5.2005
R2191 VSS.n734 VSS.n704 5.2005
R2192 VSS.n704 VSS.n117 5.2005
R2193 VSS.n736 VSS.n735 5.2005
R2194 VSS.n738 VSS.n703 5.2005
R2195 VSS.n739 VSS.n702 5.2005
R2196 VSS.n742 VSS.n741 5.2005
R2197 VSS.n214 VSS.n123 5.2005
R2198 VSS.n217 VSS.n216 5.2005
R2199 VSS.n219 VSS.n218 5.2005
R2200 VSS.n221 VSS.n213 5.2005
R2201 VSS.n222 VSS.n212 5.2005
R2202 VSS.n223 VSS.n222 5.2005
R2203 VSS.n226 VSS.n225 5.2005
R2204 VSS.n225 VSS.n224 5.2005
R2205 VSS.n227 VSS.n211 5.2005
R2206 VSS.n211 VSS.n210 5.2005
R2207 VSS.n229 VSS.n228 5.2005
R2208 VSS.n230 VSS.n229 5.2005
R2209 VSS.n209 VSS.n208 5.2005
R2210 VSS.n231 VSS.n209 5.2005
R2211 VSS.n234 VSS.n233 5.2005
R2212 VSS.n233 VSS.n232 5.2005
R2213 VSS.n235 VSS.n206 5.2005
R2214 VSS.n206 VSS.n204 5.2005
R2215 VSS.n2958 VSS.n2957 5.2005
R2216 VSS.n2959 VSS.n2958 5.2005
R2217 VSS.n2956 VSS.n207 5.2005
R2218 VSS.n207 VSS.n205 5.2005
R2219 VSS.n2955 VSS.n2954 5.2005
R2220 VSS.n2954 VSS.n2953 5.2005
R2221 VSS.n237 VSS.n236 5.2005
R2222 VSS.n2952 VSS.n237 5.2005
R2223 VSS.n2950 VSS.n2949 5.2005
R2224 VSS.n2951 VSS.n2950 5.2005
R2225 VSS.n2948 VSS.n239 5.2005
R2226 VSS.n242 VSS.n239 5.2005
R2227 VSS.n2947 VSS.n2946 5.2005
R2228 VSS.n2946 VSS.n2945 5.2005
R2229 VSS.n241 VSS.n240 5.2005
R2230 VSS.n2921 VSS.n2919 5.2005
R2231 VSS.n2922 VSS.n2918 5.2005
R2232 VSS.n2925 VSS.n2924 5.2005
R2233 VSS.n813 VSS.n812 5.2005
R2234 VSS.n812 VSS.n151 5.2005
R2235 VSS.n811 VSS.n797 5.2005
R2236 VSS.n809 VSS.n808 5.2005
R2237 VSS.n807 VSS.n798 5.2005
R2238 VSS.n806 VSS.n805 5.2005
R2239 VSS.n803 VSS.n799 5.2005
R2240 VSS.n801 VSS.n800 5.2005
R2241 VSS.n792 VSS.n791 5.2005
R2242 VSS.n792 VSS.n151 5.2005
R2243 VSS.n891 VSS.n890 5.2005
R2244 VSS.n890 VSS.n889 5.2005
R2245 VSS.n892 VSS.n790 5.2005
R2246 VSS.n793 VSS.n790 5.2005
R2247 VSS.n894 VSS.n893 5.2005
R2248 VSS.n896 VSS.n788 5.2005
R2249 VSS.n899 VSS.n898 5.2005
R2250 VSS.n898 VSS.n897 5.2005
R2251 VSS.n900 VSS.n786 5.2005
R2252 VSS.n786 VSS.n785 5.2005
R2253 VSS.n902 VSS.n901 5.2005
R2254 VSS.n903 VSS.n902 5.2005
R2255 VSS.n787 VSS.n783 5.2005
R2256 VSS.n904 VSS.n783 5.2005
R2257 VSS.n906 VSS.n784 5.2005
R2258 VSS.n906 VSS.n905 5.2005
R2259 VSS.n831 VSS.n830 5.2005
R2260 VSS.n828 VSS.n814 5.2005
R2261 VSS.n827 VSS.n826 5.2005
R2262 VSS.n825 VSS.n824 5.2005
R2263 VSS.n823 VSS.n816 5.2005
R2264 VSS.n821 VSS.n820 5.2005
R2265 VSS.n819 VSS.n818 5.2005
R2266 VSS.n155 VSS.n153 5.2005
R2267 VSS.n3056 VSS.n3055 5.2005
R2268 VSS.n3057 VSS.n3056 5.2005
R2269 VSS.n3054 VSS.n154 5.2005
R2270 VSS.n154 VSS.n152 5.2005
R2271 VSS.n3053 VSS.n3052 5.2005
R2272 VSS.n3052 VSS.n3051 5.2005
R2273 VSS.n157 VSS.n156 5.2005
R2274 VSS.n3049 VSS.n157 5.2005
R2275 VSS.n3047 VSS.n3046 5.2005
R2276 VSS.n3048 VSS.n3047 5.2005
R2277 VSS.n3045 VSS.n161 5.2005
R2278 VSS.n161 VSS.n160 5.2005
R2279 VSS.n852 VSS.n851 5.2005
R2280 VSS.n853 VSS.n845 5.2005
R2281 VSS.n855 VSS.n854 5.2005
R2282 VSS.n857 VSS.n843 5.2005
R2283 VSS.n859 VSS.n858 5.2005
R2284 VSS.n860 VSS.n842 5.2005
R2285 VSS.n862 VSS.n861 5.2005
R2286 VSS.n862 VSS.n19 5.2005
R2287 VSS.n863 VSS.n841 5.2005
R2288 VSS.n864 VSS.n863 5.2005
R2289 VSS.n867 VSS.n866 5.2005
R2290 VSS.n866 VSS.n865 5.2005
R2291 VSS.n868 VSS.n840 5.2005
R2292 VSS.n840 VSS.n839 5.2005
R2293 VSS.n870 VSS.n869 5.2005
R2294 VSS.n871 VSS.n870 5.2005
R2295 VSS.n837 VSS.n836 5.2005
R2296 VSS.n872 VSS.n837 5.2005
R2297 VSS.n875 VSS.n874 5.2005
R2298 VSS.n874 VSS.n873 5.2005
R2299 VSS.n876 VSS.n835 5.2005
R2300 VSS.n838 VSS.n835 5.2005
R2301 VSS.n878 VSS.n877 5.2005
R2302 VSS.n879 VSS.n878 5.2005
R2303 VSS.n834 VSS.n833 5.2005
R2304 VSS.n880 VSS.n834 5.2005
R2305 VSS.n883 VSS.n882 5.2005
R2306 VSS.n882 VSS.n881 5.2005
R2307 VSS.n884 VSS.n796 5.2005
R2308 VSS.n796 VSS.n794 5.2005
R2309 VSS.n886 VSS.n885 5.2005
R2310 VSS.n887 VSS.n886 5.2005
R2311 VSS.n150 VSS.n149 5.2005
R2312 VSS.n3059 VSS.n150 5.2005
R2313 VSS.n3062 VSS.n3061 5.2005
R2314 VSS.n3061 VSS.n3060 5.2005
R2315 VSS.n3063 VSS.n148 5.2005
R2316 VSS.n148 VSS.n147 5.2005
R2317 VSS.n3065 VSS.n3064 5.2005
R2318 VSS.n3066 VSS.n3065 5.2005
R2319 VSS.n146 VSS.n145 5.2005
R2320 VSS.n3067 VSS.n146 5.2005
R2321 VSS.n3070 VSS.n3069 5.2005
R2322 VSS.n3069 VSS.n3068 5.2005
R2323 VSS.n3071 VSS.n144 5.2005
R2324 VSS.n144 VSS.n143 5.2005
R2325 VSS.n3073 VSS.n3072 5.2005
R2326 VSS.n3074 VSS.n3073 5.2005
R2327 VSS.n137 VSS.n136 5.2005
R2328 VSS.n3075 VSS.n137 5.2005
R2329 VSS.n3078 VSS.n3077 5.2005
R2330 VSS.n3077 VSS.n3076 5.2005
R2331 VSS.n3079 VSS.n135 5.2005
R2332 VSS.n141 VSS.n135 5.2005
R2333 VSS.n3081 VSS.n3080 5.2005
R2334 VSS.n3083 VSS.n134 5.2005
R2335 VSS.n3084 VSS.n132 5.2005
R2336 VSS.n3087 VSS.n3086 5.2005
R2337 VSS.n3088 VSS.n131 5.2005
R2338 VSS.n131 VSS.n130 5.2005
R2339 VSS.n3090 VSS.n3089 5.2005
R2340 VSS.n3091 VSS.n3090 5.2005
R2341 VSS.n127 VSS.n125 5.2005
R2342 VSS.n3092 VSS.n127 5.2005
R2343 VSS.n3095 VSS.n3094 5.2005
R2344 VSS.n3094 VSS.n3093 5.2005
R2345 VSS.n3097 VSS.n121 5.2005
R2346 VSS.n128 VSS.n121 5.2005
R2347 VSS.n3099 VSS.n3098 5.2005
R2348 VSS.n3100 VSS.n3099 5.2005
R2349 VSS.n122 VSS.n120 5.2005
R2350 VSS.n120 VSS.n118 5.2005
R2351 VSS.n2802 VSS.n2801 5.2005
R2352 VSS.n2801 VSS.n2800 5.2005
R2353 VSS.n2804 VSS.n2803 5.2005
R2354 VSS.n2805 VSS.n2804 5.2005
R2355 VSS.n2799 VSS.n2798 5.2005
R2356 VSS.n2806 VSS.n2799 5.2005
R2357 VSS.n2809 VSS.n2808 5.2005
R2358 VSS.n2808 VSS.n2807 5.2005
R2359 VSS.n2810 VSS.n2797 5.2005
R2360 VSS.n2797 VSS.n2796 5.2005
R2361 VSS.n2812 VSS.n2811 5.2005
R2362 VSS.n2813 VSS.n2812 5.2005
R2363 VSS.n2795 VSS.n2794 5.2005
R2364 VSS.n2814 VSS.n2795 5.2005
R2365 VSS.n2817 VSS.n2816 5.2005
R2366 VSS.n2816 VSS.n2815 5.2005
R2367 VSS.n2818 VSS.n2793 5.2005
R2368 VSS.n2793 VSS.n2792 5.2005
R2369 VSS.n2820 VSS.n2819 5.2005
R2370 VSS.n2821 VSS.n2820 5.2005
R2371 VSS.n2791 VSS.n2790 5.2005
R2372 VSS.n2822 VSS.n2791 5.2005
R2373 VSS.n2825 VSS.n2824 5.2005
R2374 VSS.n2824 VSS.n2823 5.2005
R2375 VSS.n2826 VSS.n2789 5.2005
R2376 VSS.n2789 VSS.n2788 5.2005
R2377 VSS.n2828 VSS.n2827 5.2005
R2378 VSS.n2829 VSS.n2828 5.2005
R2379 VSS.n2787 VSS.n2786 5.2005
R2380 VSS.n2830 VSS.n2787 5.2005
R2381 VSS.n2833 VSS.n2832 5.2005
R2382 VSS.n2832 VSS.n2831 5.2005
R2383 VSS.n2785 VSS.n2784 5.2005
R2384 VSS.n2784 VSS.n285 5.2005
R2385 VSS.n2783 VSS.n293 5.2005
R2386 VSS.n2783 VSS.n2782 5.2005
R2387 VSS.n2777 VSS.n294 5.2005
R2388 VSS.n2781 VSS.n294 5.2005
R2389 VSS.n2779 VSS.n2778 5.2005
R2390 VSS.n2780 VSS.n2779 5.2005
R2391 VSS.n2776 VSS.n296 5.2005
R2392 VSS.n296 VSS.n295 5.2005
R2393 VSS.n2775 VSS.n2774 5.2005
R2394 VSS.n2774 VSS.n2773 5.2005
R2395 VSS.n298 VSS.n297 5.2005
R2396 VSS.n2772 VSS.n298 5.2005
R2397 VSS.n2770 VSS.n2769 5.2005
R2398 VSS.n2771 VSS.n2770 5.2005
R2399 VSS.n2768 VSS.n300 5.2005
R2400 VSS.n300 VSS.n299 5.2005
R2401 VSS.n2767 VSS.n2766 5.2005
R2402 VSS.n2766 VSS.n2765 5.2005
R2403 VSS.n302 VSS.n301 5.2005
R2404 VSS.n2764 VSS.n302 5.2005
R2405 VSS.n2762 VSS.n2761 5.2005
R2406 VSS.n2763 VSS.n2762 5.2005
R2407 VSS.n2760 VSS.n304 5.2005
R2408 VSS.n304 VSS.n303 5.2005
R2409 VSS.n2759 VSS.n2758 5.2005
R2410 VSS.n2758 VSS.n2757 5.2005
R2411 VSS.n306 VSS.n305 5.2005
R2412 VSS.n2756 VSS.n306 5.2005
R2413 VSS.n2754 VSS.n2753 5.2005
R2414 VSS.n2755 VSS.n2754 5.2005
R2415 VSS.n2752 VSS.n308 5.2005
R2416 VSS.n308 VSS.n307 5.2005
R2417 VSS.n2751 VSS.n2750 5.2005
R2418 VSS.n2750 VSS.n2749 5.2005
R2419 VSS.n310 VSS.n309 5.2005
R2420 VSS.n2748 VSS.n310 5.2005
R2421 VSS.n2532 VSS.n2531 5.2005
R2422 VSS.n2531 VSS.n355 5.2005
R2423 VSS.n2533 VSS.n2530 5.2005
R2424 VSS.n2530 VSS.n2529 5.2005
R2425 VSS.n2535 VSS.n2534 5.2005
R2426 VSS.n2536 VSS.n2535 5.2005
R2427 VSS.n2528 VSS.n2527 5.2005
R2428 VSS.n2537 VSS.n2528 5.2005
R2429 VSS.n2540 VSS.n2539 5.2005
R2430 VSS.n2539 VSS.n2538 5.2005
R2431 VSS.n2541 VSS.n2526 5.2005
R2432 VSS.n2526 VSS.n2525 5.2005
R2433 VSS.n2543 VSS.n2542 5.2005
R2434 VSS.n2544 VSS.n2543 5.2005
R2435 VSS.n2524 VSS.n2523 5.2005
R2436 VSS.n2545 VSS.n2524 5.2005
R2437 VSS.n2548 VSS.n2547 5.2005
R2438 VSS.n2547 VSS.n2546 5.2005
R2439 VSS.n2549 VSS.n2522 5.2005
R2440 VSS.n2522 VSS.n2521 5.2005
R2441 VSS.n2551 VSS.n2550 5.2005
R2442 VSS.n2552 VSS.n2551 5.2005
R2443 VSS.n2520 VSS.n2519 5.2005
R2444 VSS.n2553 VSS.n2520 5.2005
R2445 VSS.n2556 VSS.n2555 5.2005
R2446 VSS.n2555 VSS.n2554 5.2005
R2447 VSS.n2557 VSS.n2518 5.2005
R2448 VSS.n2518 VSS.n2517 5.2005
R2449 VSS.n2559 VSS.n2558 5.2005
R2450 VSS.n2560 VSS.n2559 5.2005
R2451 VSS.n2516 VSS.n2515 5.2005
R2452 VSS.n2561 VSS.n2516 5.2005
R2453 VSS.n2564 VSS.n2563 5.2005
R2454 VSS.n2563 VSS.n2562 5.2005
R2455 VSS.n2565 VSS.n438 5.2005
R2456 VSS.n438 VSS.n436 5.2005
R2457 VSS.n2567 VSS.n2566 5.2005
R2458 VSS.n2568 VSS.n2567 5.2005
R2459 VSS.n2513 VSS.n2512 5.2005
R2460 VSS.n2512 VSS.n2511 5.2005
R2461 VSS.n449 VSS.n448 5.2005
R2462 VSS.n2510 VSS.n449 5.2005
R2463 VSS.n2508 VSS.n2507 5.2005
R2464 VSS.n2509 VSS.n2508 5.2005
R2465 VSS.n2506 VSS.n451 5.2005
R2466 VSS.n451 VSS.n450 5.2005
R2467 VSS.n2505 VSS.n2504 5.2005
R2468 VSS.n2504 VSS.n2503 5.2005
R2469 VSS.n453 VSS.n452 5.2005
R2470 VSS.n2502 VSS.n453 5.2005
R2471 VSS.n2500 VSS.n2499 5.2005
R2472 VSS.n2501 VSS.n2500 5.2005
R2473 VSS.n2498 VSS.n455 5.2005
R2474 VSS.n455 VSS.n454 5.2005
R2475 VSS.n2497 VSS.n2496 5.2005
R2476 VSS.n2496 VSS.n2495 5.2005
R2477 VSS.n457 VSS.n456 5.2005
R2478 VSS.n2494 VSS.n457 5.2005
R2479 VSS.n2492 VSS.n2491 5.2005
R2480 VSS.n2493 VSS.n2492 5.2005
R2481 VSS.n2490 VSS.n459 5.2005
R2482 VSS.n459 VSS.n458 5.2005
R2483 VSS.n2489 VSS.n2488 5.2005
R2484 VSS.n2488 VSS.n2487 5.2005
R2485 VSS.n461 VSS.n460 5.2005
R2486 VSS.n2486 VSS.n461 5.2005
R2487 VSS.n2484 VSS.n2483 5.2005
R2488 VSS.n2485 VSS.n2484 5.2005
R2489 VSS.n2482 VSS.n463 5.2005
R2490 VSS.n463 VSS.n462 5.2005
R2491 VSS.n2481 VSS.n2480 5.2005
R2492 VSS.n2480 VSS.n2479 5.2005
R2493 VSS.n465 VSS.n464 5.2005
R2494 VSS.n2478 VSS.n465 5.2005
R2495 VSS.n2476 VSS.n2475 5.2005
R2496 VSS.n2477 VSS.n2476 5.2005
R2497 VSS.n2473 VSS.n2472 5.2005
R2498 VSS.n2472 VSS.n2471 5.2005
R2499 VSS.n471 VSS.n470 5.2005
R2500 VSS.n472 VSS.n471 5.2005
R2501 VSS.n2268 VSS.n2267 5.2005
R2502 VSS.n2269 VSS.n2268 5.2005
R2503 VSS.n2266 VSS.n2265 5.2005
R2504 VSS.n2270 VSS.n2266 5.2005
R2505 VSS.n2273 VSS.n2272 5.2005
R2506 VSS.n2272 VSS.n2271 5.2005
R2507 VSS.n2274 VSS.n2264 5.2005
R2508 VSS.n2264 VSS.n2263 5.2005
R2509 VSS.n2276 VSS.n2275 5.2005
R2510 VSS.n2277 VSS.n2276 5.2005
R2511 VSS.n2262 VSS.n2261 5.2005
R2512 VSS.n2278 VSS.n2262 5.2005
R2513 VSS.n2281 VSS.n2280 5.2005
R2514 VSS.n2280 VSS.n2279 5.2005
R2515 VSS.n2282 VSS.n2260 5.2005
R2516 VSS.n2260 VSS.n2259 5.2005
R2517 VSS.n2284 VSS.n2283 5.2005
R2518 VSS.n2285 VSS.n2284 5.2005
R2519 VSS.n2258 VSS.n2257 5.2005
R2520 VSS.n2286 VSS.n2258 5.2005
R2521 VSS.n2289 VSS.n2288 5.2005
R2522 VSS.n2288 VSS.n2287 5.2005
R2523 VSS.n2290 VSS.n2256 5.2005
R2524 VSS.n2256 VSS.n2255 5.2005
R2525 VSS.n2292 VSS.n2291 5.2005
R2526 VSS.n2293 VSS.n2292 5.2005
R2527 VSS.n2254 VSS.n2253 5.2005
R2528 VSS.n2294 VSS.n2254 5.2005
R2529 VSS.n2297 VSS.n2296 5.2005
R2530 VSS.n2296 VSS.n2295 5.2005
R2531 VSS.n2298 VSS.n559 5.2005
R2532 VSS.n559 VSS.n557 5.2005
R2533 VSS.n2300 VSS.n2299 5.2005
R2534 VSS.n2301 VSS.n2300 5.2005
R2535 VSS.n2251 VSS.n2250 5.2005
R2536 VSS.n2250 VSS.n2249 5.2005
R2537 VSS.n570 VSS.n569 5.2005
R2538 VSS.n2248 VSS.n570 5.2005
R2539 VSS.n2246 VSS.n2245 5.2005
R2540 VSS.n2247 VSS.n2246 5.2005
R2541 VSS.n2244 VSS.n572 5.2005
R2542 VSS.n572 VSS.n571 5.2005
R2543 VSS.n2243 VSS.n2242 5.2005
R2544 VSS.n2242 VSS.n2241 5.2005
R2545 VSS.n574 VSS.n573 5.2005
R2546 VSS.n2240 VSS.n574 5.2005
R2547 VSS.n2238 VSS.n2237 5.2005
R2548 VSS.n2239 VSS.n2238 5.2005
R2549 VSS.n2236 VSS.n576 5.2005
R2550 VSS.n576 VSS.n575 5.2005
R2551 VSS.n2235 VSS.n2234 5.2005
R2552 VSS.n2234 VSS.n2233 5.2005
R2553 VSS.n578 VSS.n577 5.2005
R2554 VSS.n2232 VSS.n578 5.2005
R2555 VSS.n2230 VSS.n2229 5.2005
R2556 VSS.n2231 VSS.n2230 5.2005
R2557 VSS.n2228 VSS.n580 5.2005
R2558 VSS.n580 VSS.n579 5.2005
R2559 VSS.n2227 VSS.n2226 5.2005
R2560 VSS.n2226 VSS.n2225 5.2005
R2561 VSS.n582 VSS.n581 5.2005
R2562 VSS.n2224 VSS.n582 5.2005
R2563 VSS.n2222 VSS.n2221 5.2005
R2564 VSS.n2223 VSS.n2222 5.2005
R2565 VSS.n2220 VSS.n584 5.2005
R2566 VSS.n584 VSS.n583 5.2005
R2567 VSS.n2219 VSS.n2218 5.2005
R2568 VSS.n2218 VSS.n2217 5.2005
R2569 VSS.n586 VSS.n585 5.2005
R2570 VSS.n2214 VSS.n586 5.2005
R2571 VSS.n2212 VSS.n2211 5.2005
R2572 VSS.n2213 VSS.n2212 5.2005
R2573 VSS.n2129 VSS.n2128 5.2005
R2574 VSS.n2129 VSS.n554 5.2005
R2575 VSS.n2127 VSS.n1771 5.2005
R2576 VSS.n1815 VSS.n1771 5.2005
R2577 VSS.n2126 VSS.n2125 5.2005
R2578 VSS.n2125 VSS.n2124 5.2005
R2579 VSS.n1814 VSS.n1813 5.2005
R2580 VSS.n2123 VSS.n1814 5.2005
R2581 VSS.n2121 VSS.n2120 5.2005
R2582 VSS.n2122 VSS.n2121 5.2005
R2583 VSS.n2119 VSS.n1817 5.2005
R2584 VSS.n1817 VSS.n1816 5.2005
R2585 VSS.n2118 VSS.n2117 5.2005
R2586 VSS.n2117 VSS.n2116 5.2005
R2587 VSS.n1819 VSS.n1818 5.2005
R2588 VSS.n2115 VSS.n1819 5.2005
R2589 VSS.n2113 VSS.n2112 5.2005
R2590 VSS.n2114 VSS.n2113 5.2005
R2591 VSS.n2111 VSS.n1821 5.2005
R2592 VSS.n1821 VSS.n1820 5.2005
R2593 VSS.n2110 VSS.n2109 5.2005
R2594 VSS.n2109 VSS.n2108 5.2005
R2595 VSS.n1823 VSS.n1822 5.2005
R2596 VSS.n2107 VSS.n1823 5.2005
R2597 VSS.n2105 VSS.n2104 5.2005
R2598 VSS.n2106 VSS.n2105 5.2005
R2599 VSS.n2103 VSS.n1825 5.2005
R2600 VSS.n1825 VSS.n1824 5.2005
R2601 VSS.n2102 VSS.n2101 5.2005
R2602 VSS.n2101 VSS.n2100 5.2005
R2603 VSS.n1827 VSS.n1826 5.2005
R2604 VSS.n2099 VSS.n1827 5.2005
R2605 VSS.n2097 VSS.n2096 5.2005
R2606 VSS.n2098 VSS.n2097 5.2005
R2607 VSS.n2095 VSS.n1829 5.2005
R2608 VSS.n1829 VSS.n1828 5.2005
R2609 VSS.n2094 VSS.n2093 5.2005
R2610 VSS.n2093 VSS.n2092 5.2005
R2611 VSS.n2051 VSS.n1832 5.2005
R2612 VSS.n2051 VSS.n2050 5.2005
R2613 VSS.n1835 VSS.n1831 5.2005
R2614 VSS.n2049 VSS.n1831 5.2005
R2615 VSS.n2047 VSS.n2046 5.2005
R2616 VSS.n2048 VSS.n2047 5.2005
R2617 VSS.n2045 VSS.n1834 5.2005
R2618 VSS.n1834 VSS.n1833 5.2005
R2619 VSS.n2044 VSS.n2043 5.2005
R2620 VSS.n2043 VSS.n2042 5.2005
R2621 VSS.n1837 VSS.n1836 5.2005
R2622 VSS.n2041 VSS.n1837 5.2005
R2623 VSS.n2039 VSS.n2038 5.2005
R2624 VSS.n2040 VSS.n2039 5.2005
R2625 VSS.n2037 VSS.n1839 5.2005
R2626 VSS.n1839 VSS.n1838 5.2005
R2627 VSS.n2036 VSS.n2035 5.2005
R2628 VSS.n2035 VSS.n2034 5.2005
R2629 VSS.n1841 VSS.n1840 5.2005
R2630 VSS.n2033 VSS.n1841 5.2005
R2631 VSS.n2031 VSS.n2030 5.2005
R2632 VSS.n2032 VSS.n2031 5.2005
R2633 VSS.n2029 VSS.n1843 5.2005
R2634 VSS.n1843 VSS.n1842 5.2005
R2635 VSS.n2028 VSS.n2027 5.2005
R2636 VSS.n2027 VSS.n2026 5.2005
R2637 VSS.n1845 VSS.n1844 5.2005
R2638 VSS.n2025 VSS.n1845 5.2005
R2639 VSS.n2023 VSS.n2022 5.2005
R2640 VSS.n2024 VSS.n2023 5.2005
R2641 VSS.n2021 VSS.n1847 5.2005
R2642 VSS.n1847 VSS.n1846 5.2005
R2643 VSS.n2020 VSS.n2019 5.2005
R2644 VSS.n2019 VSS.n2018 5.2005
R2645 VSS.n1849 VSS.n1848 5.2005
R2646 VSS.n2017 VSS.n1849 5.2005
R2647 VSS.n2015 VSS.n2014 5.2005
R2648 VSS.n2016 VSS.n2015 5.2005
R2649 VSS.n2012 VSS.n2011 5.2005
R2650 VSS.n2011 VSS.n434 5.2005
R2651 VSS.n2010 VSS.n1892 5.2005
R2652 VSS.n2010 VSS.n2009 5.2005
R2653 VSS.n1896 VSS.n1893 5.2005
R2654 VSS.n2008 VSS.n1893 5.2005
R2655 VSS.n2006 VSS.n2005 5.2005
R2656 VSS.n2007 VSS.n2006 5.2005
R2657 VSS.n2004 VSS.n1895 5.2005
R2658 VSS.n1895 VSS.n1894 5.2005
R2659 VSS.n2003 VSS.n2002 5.2005
R2660 VSS.n2002 VSS.n2001 5.2005
R2661 VSS.n1898 VSS.n1897 5.2005
R2662 VSS.n2000 VSS.n1898 5.2005
R2663 VSS.n1998 VSS.n1997 5.2005
R2664 VSS.n1999 VSS.n1998 5.2005
R2665 VSS.n1996 VSS.n1900 5.2005
R2666 VSS.n1900 VSS.n1899 5.2005
R2667 VSS.n1995 VSS.n1994 5.2005
R2668 VSS.n1994 VSS.n1993 5.2005
R2669 VSS.n1902 VSS.n1901 5.2005
R2670 VSS.n1992 VSS.n1902 5.2005
R2671 VSS.n1990 VSS.n1989 5.2005
R2672 VSS.n1991 VSS.n1990 5.2005
R2673 VSS.n1988 VSS.n1904 5.2005
R2674 VSS.n1904 VSS.n1903 5.2005
R2675 VSS.n1987 VSS.n1986 5.2005
R2676 VSS.n1986 VSS.n1985 5.2005
R2677 VSS.n1906 VSS.n1905 5.2005
R2678 VSS.n1984 VSS.n1906 5.2005
R2679 VSS.n1982 VSS.n1981 5.2005
R2680 VSS.n1983 VSS.n1982 5.2005
R2681 VSS.n1980 VSS.n1908 5.2005
R2682 VSS.n1908 VSS.n1907 5.2005
R2683 VSS.n1979 VSS.n1978 5.2005
R2684 VSS.n1978 VSS.n1977 5.2005
R2685 VSS.n1975 VSS.n1909 5.2005
R2686 VSS.n1976 VSS.n1975 5.2005
R2687 VSS.n1973 VSS.n1972 5.2005
R2688 VSS.n1973 VSS.n312 5.2005
R2689 VSS.n1971 VSS.n1911 5.2005
R2690 VSS.n1954 VSS.n1911 5.2005
R2691 VSS.n1970 VSS.n1969 5.2005
R2692 VSS.n1969 VSS.n1968 5.2005
R2693 VSS.n1953 VSS.n1952 5.2005
R2694 VSS.n1967 VSS.n1953 5.2005
R2695 VSS.n1965 VSS.n1964 5.2005
R2696 VSS.n1966 VSS.n1965 5.2005
R2697 VSS.n1963 VSS.n1956 5.2005
R2698 VSS.n1956 VSS.n1955 5.2005
R2699 VSS.n1962 VSS.n1961 5.2005
R2700 VSS.n1961 VSS.n1960 5.2005
R2701 VSS.n1958 VSS.n1957 5.2005
R2702 VSS.n1959 VSS.n1958 5.2005
R2703 VSS.n85 VSS.n83 5.2005
R2704 VSS.n83 VSS.n79 5.2005
R2705 VSS.n3156 VSS.n3155 5.2005
R2706 VSS.n3157 VSS.n3156 5.2005
R2707 VSS.n3154 VSS.n84 5.2005
R2708 VSS.n88 VSS.n84 5.2005
R2709 VSS.n3153 VSS.n3152 5.2005
R2710 VSS.n3152 VSS.n3151 5.2005
R2711 VSS.n87 VSS.n86 5.2005
R2712 VSS.n3150 VSS.n87 5.2005
R2713 VSS.n3148 VSS.n3147 5.2005
R2714 VSS.n3149 VSS.n3148 5.2005
R2715 VSS.n3146 VSS.n90 5.2005
R2716 VSS.n90 VSS.n89 5.2005
R2717 VSS.n3145 VSS.n3144 5.2005
R2718 VSS.n3144 VSS.n3143 5.2005
R2719 VSS.n92 VSS.n91 5.2005
R2720 VSS.n3142 VSS.n92 5.2005
R2721 VSS.n3140 VSS.n3139 5.2005
R2722 VSS.n3141 VSS.n3140 5.2005
R2723 VSS.n3138 VSS.n94 5.2005
R2724 VSS.n94 VSS.n93 5.2005
R2725 VSS.n3136 VSS.n3135 5.2005
R2726 VSS.n3135 VSS.n3134 5.2005
R2727 VSS.n98 VSS.n96 5.2005
R2728 VSS.n3133 VSS.n98 5.2005
R2729 VSS.n3131 VSS.n3130 5.2005
R2730 VSS.n3132 VSS.n3131 5.2005
R2731 VSS.n3129 VSS.n101 5.2005
R2732 VSS.n101 VSS.n100 5.2005
R2733 VSS.n3128 VSS.n3127 5.2005
R2734 VSS.n3127 VSS.n3126 5.2005
R2735 VSS.n103 VSS.n102 5.2005
R2736 VSS.n3125 VSS.n103 5.2005
R2737 VSS.n3123 VSS.n3122 5.2005
R2738 VSS.n3124 VSS.n3123 5.2005
R2739 VSS.n3121 VSS.n105 5.2005
R2740 VSS.n105 VSS.n104 5.2005
R2741 VSS.n3120 VSS.n3119 5.2005
R2742 VSS.n3119 VSS.n3118 5.2005
R2743 VSS.n107 VSS.n106 5.2005
R2744 VSS.n3117 VSS.n107 5.2005
R2745 VSS.n3115 VSS.n3114 5.2005
R2746 VSS.n3116 VSS.n3115 5.2005
R2747 VSS.n3113 VSS.n108 5.2005
R2748 VSS.n111 VSS.n108 5.2005
R2749 VSS.n3112 VSS.n3111 5.2005
R2750 VSS.n3111 VSS.n3110 5.2005
R2751 VSS.n110 VSS.n109 5.2005
R2752 VSS.n3109 VSS.n110 5.2005
R2753 VSS.n3107 VSS.n3106 5.2005
R2754 VSS.n3108 VSS.n3107 5.2005
R2755 VSS.n3105 VSS.n113 5.2005
R2756 VSS.n113 VSS.n112 5.2005
R2757 VSS.n3104 VSS.n3103 5.2005
R2758 VSS.n3103 VSS.n3102 5.2005
R2759 VSS.n115 VSS.n114 5.2005
R2760 VSS.n116 VSS.n115 5.2005
R2761 VSS.n745 VSS.n744 5.2005
R2762 VSS.n744 VSS.n743 5.2005
R2763 VSS.n748 VSS.n747 5.2005
R2764 VSS.n749 VSS.n748 5.2005
R2765 VSS.n699 VSS.n698 5.2005
R2766 VSS.n750 VSS.n699 5.2005
R2767 VSS.n753 VSS.n752 5.2005
R2768 VSS.n752 VSS.n751 5.2005
R2769 VSS.n754 VSS.n697 5.2005
R2770 VSS.n697 VSS.n70 5.2005
R2771 VSS.n756 VSS.n755 5.2005
R2772 VSS.n758 VSS.n696 5.2005
R2773 VSS.n759 VSS.n695 5.2005
R2774 VSS.n759 VSS.n81 5.2005
R2775 VSS.n762 VSS.n761 5.2005
R2776 VSS.n763 VSS.n694 5.2005
R2777 VSS.n765 VSS.n764 5.2005
R2778 VSS.n765 VSS.n81 5.2005
R2779 VSS.n766 VSS.n693 5.2005
R2780 VSS.n769 VSS.n768 5.2005
R2781 VSS.n770 VSS.n692 5.2005
R2782 VSS.n692 VSS.n80 5.2005
R2783 VSS.n772 VSS.n771 5.2005
R2784 VSS.n774 VSS.n691 5.2005
R2785 VSS.n777 VSS.n776 5.2005
R2786 VSS.n778 VSS.n690 5.2005
R2787 VSS.n780 VSS.n779 5.2005
R2788 VSS.n782 VSS.n689 5.2005
R2789 VSS.n910 VSS.n909 5.2005
R2790 VSS.n911 VSS.n687 5.2005
R2791 VSS.n913 VSS.n912 5.2005
R2792 VSS.n915 VSS.n686 5.2005
R2793 VSS.n918 VSS.n917 5.2005
R2794 VSS.n919 VSS.n685 5.2005
R2795 VSS.n921 VSS.n920 5.2005
R2796 VSS.n923 VSS.n684 5.2005
R2797 VSS.n926 VSS.n925 5.2005
R2798 VSS.n927 VSS.n683 5.2005
R2799 VSS.n929 VSS.n928 5.2005
R2800 VSS.n931 VSS.n682 5.2005
R2801 VSS.n934 VSS.n933 5.2005
R2802 VSS.n935 VSS.n681 5.2005
R2803 VSS.n937 VSS.n936 5.2005
R2804 VSS.n939 VSS.n680 5.2005
R2805 VSS.n942 VSS.n941 5.2005
R2806 VSS.n943 VSS.n679 5.2005
R2807 VSS.n945 VSS.n944 5.2005
R2808 VSS.n945 VSS.n80 5.2005
R2809 VSS.n1661 VSS.n1660 5.2005
R2810 VSS.n1663 VSS.n1662 5.2005
R2811 VSS.n1665 VSS.n1664 5.2005
R2812 VSS.n1667 VSS.n1666 5.2005
R2813 VSS.n1669 VSS.n1668 5.2005
R2814 VSS.n1671 VSS.n1670 5.2005
R2815 VSS.n1673 VSS.n1672 5.2005
R2816 VSS.n1675 VSS.n1674 5.2005
R2817 VSS.n1677 VSS.n1676 5.2005
R2818 VSS.n1679 VSS.n1678 5.2005
R2819 VSS.n1681 VSS.n1680 5.2005
R2820 VSS.n1683 VSS.n1682 5.2005
R2821 VSS.n1685 VSS.n1684 5.2005
R2822 VSS.n1686 VSS.n1070 5.2005
R2823 VSS.n1688 VSS.n1687 5.2005
R2824 VSS.n1060 VSS.n1058 5.2005
R2825 VSS.n1692 VSS.n1691 5.2005
R2826 VSS.n1691 VSS.n1690 5.2005
R2827 VSS.n1287 VSS.n1263 5.2005
R2828 VSS.n1267 VSS.n1263 5.2005
R2829 VSS.n1286 VSS.n1285 5.2005
R2830 VSS.n1285 VSS.n1284 5.2005
R2831 VSS.n1266 VSS.n1265 5.2005
R2832 VSS.n1283 VSS.n1266 5.2005
R2833 VSS.n1281 VSS.n1280 5.2005
R2834 VSS.n1282 VSS.n1281 5.2005
R2835 VSS.n1279 VSS.n1269 5.2005
R2836 VSS.n1269 VSS.n1268 5.2005
R2837 VSS.n1278 VSS.n1277 5.2005
R2838 VSS.n1277 VSS.n1276 5.2005
R2839 VSS.n1274 VSS.n1270 5.2005
R2840 VSS.n1275 VSS.n1274 5.2005
R2841 VSS.n1273 VSS.n1272 5.2005
R2842 VSS.n1273 VSS.n1076 5.2005
R2843 VSS.n1271 VSS.n1059 5.2005
R2844 VSS.n1061 VSS.n1059 5.2005
R2845 VSS.n1659 VSS.n1658 5.2005
R2846 VSS.n1659 VSS.n1061 5.2005
R2847 VSS.n1249 VSS.n1248 5.2005
R2848 VSS.n1251 VSS.n1250 5.2005
R2849 VSS.n1244 VSS.n1241 5.2005
R2850 VSS.n1246 VSS.n1245 5.2005
R2851 VSS.n1245 VSS.n1210 5.2005
R2852 VSS.n1202 VSS.n1201 5.2005
R2853 VSS.n1199 VSS.n1165 5.2005
R2854 VSS.n1199 VSS.n1161 5.2005
R2855 VSS.n1198 VSS.n1197 5.2005
R2856 VSS.n1196 VSS.n1195 5.2005
R2857 VSS.n1194 VSS.n1167 5.2005
R2858 VSS.n1192 VSS.n1191 5.2005
R2859 VSS.n1190 VSS.n1168 5.2005
R2860 VSS.n1189 VSS.n1188 5.2005
R2861 VSS.n1186 VSS.n1169 5.2005
R2862 VSS.n1184 VSS.n1183 5.2005
R2863 VSS.n1182 VSS.n1170 5.2005
R2864 VSS.n1181 VSS.n1180 5.2005
R2865 VSS.n1178 VSS.n1171 5.2005
R2866 VSS.n1176 VSS.n1175 5.2005
R2867 VSS.n1174 VSS.n1173 5.2005
R2868 VSS.n1159 VSS.n1156 5.2005
R2869 VSS.n1312 VSS.n1311 5.2005
R2870 VSS.n1314 VSS.n1313 5.2005
R2871 VSS.n1316 VSS.n1315 5.2005
R2872 VSS.n1318 VSS.n1317 5.2005
R2873 VSS.n1320 VSS.n1319 5.2005
R2874 VSS.n1322 VSS.n1321 5.2005
R2875 VSS.n1324 VSS.n1323 5.2005
R2876 VSS.n1326 VSS.n1325 5.2005
R2877 VSS.n1328 VSS.n1327 5.2005
R2878 VSS.n1330 VSS.n1329 5.2005
R2879 VSS.n1332 VSS.n1331 5.2005
R2880 VSS.n1334 VSS.n1333 5.2005
R2881 VSS.n1336 VSS.n1335 5.2005
R2882 VSS.n1338 VSS.n1337 5.2005
R2883 VSS.n1340 VSS.n1339 5.2005
R2884 VSS.n1341 VSS.n1237 5.2005
R2885 VSS.n1343 VSS.n1342 5.2005
R2886 VSS.n1344 VSS.n1343 5.2005
R2887 VSS.n1307 VSS.n1291 5.2005
R2888 VSS.n1291 VSS.n1290 5.2005
R2889 VSS.n1309 VSS.n1308 5.2005
R2890 VSS.n1309 VSS.n1228 5.2005
R2891 VSS.n1260 VSS.n1227 5.2005
R2892 VSS.n1345 VSS.n1227 5.2005
R2893 VSS.n1259 VSS.n1258 5.2005
R2894 VSS.n1258 VSS.n1222 5.2005
R2895 VSS.n1257 VSS.n1221 5.2005
R2896 VSS.n1351 VSS.n1221 5.2005
R2897 VSS.n1256 VSS.n1220 5.2005
R2898 VSS.n1361 VSS.n1220 5.2005
R2899 VSS.n1255 VSS.n1219 5.2005
R2900 VSS.n1362 VSS.n1219 5.2005
R2901 VSS.n1254 VSS.n1253 5.2005
R2902 VSS.n1253 VSS.n1252 5.2005
R2903 VSS.n1240 VSS.n1209 5.2005
R2904 VSS.n1367 VSS.n1209 5.2005
R2905 VSS.n1239 VSS.n1208 5.2005
R2906 VSS.n1368 VSS.n1208 5.2005
R2907 VSS.n1238 VSS.n1207 5.2005
R2908 VSS.n1369 VSS.n1207 5.2005
R2909 VSS.n1160 VSS.n1158 5.2005
R2910 VSS.n1162 VSS.n1160 5.2005
R2911 VSS.n1377 VSS.n1376 5.2005
R2912 VSS.n1376 VSS.n1375 5.2005
R2913 VSS.n1374 VSS.n1373 5.2005
R2914 VSS.n1375 VSS.n1374 5.2005
R2915 VSS.n1372 VSS.n1164 5.2005
R2916 VSS.n1164 VSS.n1162 5.2005
R2917 VSS.n1371 VSS.n1370 5.2005
R2918 VSS.n1370 VSS.n1369 5.2005
R2919 VSS.n1206 VSS.n1205 5.2005
R2920 VSS.n1368 VSS.n1206 5.2005
R2921 VSS.n1367 VSS.n1366 5.2005
R2922 VSS.n1252 VSS.n1211 5.2005
R2923 VSS.n1364 VSS.n1363 5.2005
R2924 VSS.n1363 VSS.n1362 5.2005
R2925 VSS.n1224 VSS.n1217 5.2005
R2926 VSS.n1361 VSS.n1217 5.2005
R2927 VSS.n1350 VSS.n1349 5.2005
R2928 VSS.n1351 VSS.n1350 5.2005
R2929 VSS.n1348 VSS.n1223 5.2005
R2930 VSS.n1223 VSS.n1222 5.2005
R2931 VSS.n1347 VSS.n1346 5.2005
R2932 VSS.n1346 VSS.n1345 5.2005
R2933 VSS.n1264 VSS.n1262 5.2005
R2934 VSS.n1262 VSS.n1228 5.2005
R2935 VSS.n1289 VSS.n1288 5.2005
R2936 VSS.n1290 VSS.n1289 5.2005
R2937 VSS.n1656 VSS.n1655 5.2005
R2938 VSS.n1655 VSS.n1654 5.2005
R2939 VSS.n1074 VSS.n1073 5.2005
R2940 VSS.n1075 VSS.n1074 5.2005
R2941 VSS.n1298 VSS.n1297 5.2005
R2942 VSS.n1297 VSS.n1296 5.2005
R2943 VSS.n1299 VSS.n1295 5.2005
R2944 VSS.n1295 VSS.n1294 5.2005
R2945 VSS.n1301 VSS.n1300 5.2005
R2946 VSS.n1302 VSS.n1301 5.2005
R2947 VSS.n1293 VSS.n1292 5.2005
R2948 VSS.n1303 VSS.n1293 5.2005
R2949 VSS.n1306 VSS.n1305 5.2005
R2950 VSS.n1305 VSS.n1304 5.2005
R2951 VSS.n1657 VSS.n1072 5.2005
R2952 VSS.n1497 VSS.n1496 5.2005
R2953 VSS.n1499 VSS.n1498 5.2005
R2954 VSS.n1501 VSS.n1500 5.2005
R2955 VSS.n1502 VSS.n1453 5.2005
R2956 VSS.n1504 VSS.n1503 5.2005
R2957 VSS.n1505 VSS.n1504 5.2005
R2958 VSS.n1495 VSS.n1452 5.2005
R2959 VSS.n1452 VSS.n1451 5.2005
R2960 VSS.n1494 VSS.n1493 5.2005
R2961 VSS.n1493 VSS.n1492 5.2005
R2962 VSS.n1455 VSS.n1454 5.2005
R2963 VSS.n1491 VSS.n1455 5.2005
R2964 VSS.n1489 VSS.n1488 5.2005
R2965 VSS.n1490 VSS.n1489 5.2005
R2966 VSS.n1487 VSS.n1457 5.2005
R2967 VSS.n1457 VSS.n1456 5.2005
R2968 VSS.n1486 VSS.n1485 5.2005
R2969 VSS.n1485 VSS.n1443 5.2005
R2970 VSS.n1484 VSS.n1483 5.2005
R2971 VSS.n1484 VSS.n1442 5.2005
R2972 VSS.n1482 VSS.n1458 5.2005
R2973 VSS.n1478 VSS.n1458 5.2005
R2974 VSS.n1481 VSS.n1480 5.2005
R2975 VSS.n1480 VSS.n1479 5.2005
R2976 VSS.n1460 VSS.n1459 5.2005
R2977 VSS.n1477 VSS.n1460 5.2005
R2978 VSS.n1475 VSS.n1474 5.2005
R2979 VSS.n1476 VSS.n1475 5.2005
R2980 VSS.n1473 VSS.n1462 5.2005
R2981 VSS.n1462 VSS.n1461 5.2005
R2982 VSS.n1472 VSS.n1471 5.2005
R2983 VSS.n1471 VSS.n590 5.2005
R2984 VSS.n1470 VSS.n1468 5.2005
R2985 VSS.n1467 VSS.n1416 5.2005
R2986 VSS.n1466 VSS.n1415 5.2005
R2987 VSS.n1465 VSS.n1464 5.2005
R2988 VSS.n2194 VSS.n2193 5.2005
R2989 VSS.n2195 VSS.n2191 5.2005
R2990 VSS.n2197 VSS.n2196 5.2005
R2991 VSS.n2199 VSS.n2189 5.2005
R2992 VSS.n2201 VSS.n2200 5.2005
R2993 VSS.n2202 VSS.n2188 5.2005
R2994 VSS.n2204 VSS.n2203 5.2005
R2995 VSS.n2206 VSS.n2187 5.2005
R2996 VSS.n2208 VSS.n2207 5.2005
R2997 VSS.n2185 VSS.n596 5.2005
R2998 VSS.n2184 VSS.n2183 5.2005
R2999 VSS.n2182 VSS.n2181 5.2005
R3000 VSS.n2180 VSS.n599 5.2005
R3001 VSS.n2180 VSS.n589 5.2005
R3002 VSS.n2179 VSS.n2178 5.2005
R3003 VSS.n2177 VSS.n2176 5.2005
R3004 VSS.n2175 VSS.n601 5.2005
R3005 VSS.n616 VSS.n602 5.2005
R3006 VSS.n2171 VSS.n2170 5.2005
R3007 VSS.n2172 VSS.n2171 5.2005
R3008 VSS.n2169 VSS.n605 5.2005
R3009 VSS.n605 VSS.n587 5.2005
R3010 VSS.n2168 VSS.n2167 5.2005
R3011 VSS.n2167 VSS.n588 5.2005
R3012 VSS.n2166 VSS.n606 5.2005
R3013 VSS.n2166 VSS.n2165 5.2005
R3014 VSS.n610 VSS.n607 5.2005
R3015 VSS.n2164 VSS.n607 5.2005
R3016 VSS.n2162 VSS.n2161 5.2005
R3017 VSS.n2163 VSS.n2162 5.2005
R3018 VSS.n2160 VSS.n609 5.2005
R3019 VSS.n609 VSS.n608 5.2005
R3020 VSS.n2159 VSS.n2158 5.2005
R3021 VSS.n2158 VSS.n2157 5.2005
R3022 VSS.n612 VSS.n611 5.2005
R3023 VSS.n2156 VSS.n612 5.2005
R3024 VSS.n2150 VSS.n1761 5.2005
R3025 VSS.n2150 VSS.n2149 5.2005
R3026 VSS.n1764 VSS.n1760 5.2005
R3027 VSS.n2148 VSS.n1760 5.2005
R3028 VSS.n2146 VSS.n2145 5.2005
R3029 VSS.n2147 VSS.n2146 5.2005
R3030 VSS.n2144 VSS.n1763 5.2005
R3031 VSS.n1763 VSS.n1762 5.2005
R3032 VSS.n2143 VSS.n2142 5.2005
R3033 VSS.n2142 VSS.n2141 5.2005
R3034 VSS.n1766 VSS.n1765 5.2005
R3035 VSS.n2140 VSS.n1766 5.2005
R3036 VSS.n2138 VSS.n2137 5.2005
R3037 VSS.n2139 VSS.n2138 5.2005
R3038 VSS.n2136 VSS.n1768 5.2005
R3039 VSS.n1768 VSS.n1767 5.2005
R3040 VSS.n2135 VSS.n2134 5.2005
R3041 VSS.n2134 VSS.n2133 5.2005
R3042 VSS.n2131 VSS.n1769 5.2005
R3043 VSS.n2132 VSS.n2131 5.2005
R3044 VSS.n1554 VSS.n1553 5.2005
R3045 VSS.n1555 VSS.n1554 5.2005
R3046 VSS.n1552 VSS.n1447 5.2005
R3047 VSS.n1447 VSS.n1446 5.2005
R3048 VSS.n1551 VSS.n1550 5.2005
R3049 VSS.n1550 VSS.n1549 5.2005
R3050 VSS.n1450 VSS.n1449 5.2005
R3051 VSS.n1548 VSS.n1450 5.2005
R3052 VSS.n1546 VSS.n1545 5.2005
R3053 VSS.n1547 VSS.n1546 5.2005
R3054 VSS.n1544 VSS.n1508 5.2005
R3055 VSS.n1508 VSS.n1507 5.2005
R3056 VSS.n1543 VSS.n1542 5.2005
R3057 VSS.n1542 VSS.n1541 5.2005
R3058 VSS.n1510 VSS.n1509 5.2005
R3059 VSS.n1540 VSS.n1510 5.2005
R3060 VSS.n1538 VSS.n1537 5.2005
R3061 VSS.n1539 VSS.n1538 5.2005
R3062 VSS.n1535 VSS.n1512 5.2005
R3063 VSS.n1512 VSS.n1511 5.2005
R3064 VSS.n1534 VSS.n1533 5.2005
R3065 VSS.n1533 VSS.n1532 5.2005
R3066 VSS.n1515 VSS.n1514 5.2005
R3067 VSS.n1531 VSS.n1515 5.2005
R3068 VSS.n1529 VSS.n1528 5.2005
R3069 VSS.n1530 VSS.n1529 5.2005
R3070 VSS.n1527 VSS.n1517 5.2005
R3071 VSS.n1517 VSS.n1516 5.2005
R3072 VSS.n1526 VSS.n1525 5.2005
R3073 VSS.n1525 VSS.n1524 5.2005
R3074 VSS.n1519 VSS.n1518 5.2005
R3075 VSS.n1523 VSS.n1519 5.2005
R3076 VSS.n1521 VSS.n1520 5.2005
R3077 VSS.n1522 VSS.n1521 5.2005
R3078 VSS.n532 VSS.n531 5.2005
R3079 VSS.n533 VSS.n532 5.2005
R3080 VSS.n2342 VSS.n2341 5.2005
R3081 VSS.n2341 VSS.n2340 5.2005
R3082 VSS.n2345 VSS.n2344 5.2005
R3083 VSS.n2346 VSS.n2345 5.2005
R3084 VSS.n527 VSS.n526 5.2005
R3085 VSS.n2347 VSS.n527 5.2005
R3086 VSS.n2350 VSS.n2349 5.2005
R3087 VSS.n2349 VSS.n2348 5.2005
R3088 VSS.n2351 VSS.n525 5.2005
R3089 VSS.n525 VSS.n524 5.2005
R3090 VSS.n2353 VSS.n2352 5.2005
R3091 VSS.n2354 VSS.n2353 5.2005
R3092 VSS.n523 VSS.n522 5.2005
R3093 VSS.n2355 VSS.n523 5.2005
R3094 VSS.n2358 VSS.n2357 5.2005
R3095 VSS.n2357 VSS.n2356 5.2005
R3096 VSS.n2359 VSS.n521 5.2005
R3097 VSS.n521 VSS.n520 5.2005
R3098 VSS.n2363 VSS.n2362 5.2005
R3099 VSS.n2364 VSS.n2363 5.2005
R3100 VSS.n519 VSS.n518 5.2005
R3101 VSS.n2365 VSS.n519 5.2005
R3102 VSS.n2368 VSS.n2367 5.2005
R3103 VSS.n2367 VSS.n2366 5.2005
R3104 VSS.n2369 VSS.n517 5.2005
R3105 VSS.n517 VSS.n516 5.2005
R3106 VSS.n2371 VSS.n2370 5.2005
R3107 VSS.n2372 VSS.n2371 5.2005
R3108 VSS.n515 VSS.n514 5.2005
R3109 VSS.n2373 VSS.n515 5.2005
R3110 VSS.n2376 VSS.n2375 5.2005
R3111 VSS.n2375 VSS.n2374 5.2005
R3112 VSS.n2377 VSS.n513 5.2005
R3113 VSS.n513 VSS.n512 5.2005
R3114 VSS.n2379 VSS.n2378 5.2005
R3115 VSS.n2380 VSS.n2379 5.2005
R3116 VSS.n511 VSS.n510 5.2005
R3117 VSS.n2381 VSS.n511 5.2005
R3118 VSS.n2384 VSS.n2383 5.2005
R3119 VSS.n2383 VSS.n2382 5.2005
R3120 VSS.n2435 VSS.n2434 5.2005
R3121 VSS.n2436 VSS.n2435 5.2005
R3122 VSS.n2433 VSS.n499 5.2005
R3123 VSS.n499 VSS.n497 5.2005
R3124 VSS.n2432 VSS.n2431 5.2005
R3125 VSS.n2431 VSS.n2430 5.2005
R3126 VSS.n2387 VSS.n2386 5.2005
R3127 VSS.n2429 VSS.n2387 5.2005
R3128 VSS.n2427 VSS.n2426 5.2005
R3129 VSS.n2428 VSS.n2427 5.2005
R3130 VSS.n2425 VSS.n2389 5.2005
R3131 VSS.n2389 VSS.n2388 5.2005
R3132 VSS.n2424 VSS.n2423 5.2005
R3133 VSS.n2423 VSS.n2422 5.2005
R3134 VSS.n2391 VSS.n2390 5.2005
R3135 VSS.n2421 VSS.n2391 5.2005
R3136 VSS.n2419 VSS.n2418 5.2005
R3137 VSS.n2420 VSS.n2419 5.2005
R3138 VSS.n2416 VSS.n2393 5.2005
R3139 VSS.n2393 VSS.n2392 5.2005
R3140 VSS.n2415 VSS.n2414 5.2005
R3141 VSS.n2414 VSS.n2413 5.2005
R3142 VSS.n2396 VSS.n2395 5.2005
R3143 VSS.n2412 VSS.n2396 5.2005
R3144 VSS.n2410 VSS.n2409 5.2005
R3145 VSS.n2411 VSS.n2410 5.2005
R3146 VSS.n2408 VSS.n2398 5.2005
R3147 VSS.n2398 VSS.n2397 5.2005
R3148 VSS.n2407 VSS.n2406 5.2005
R3149 VSS.n2406 VSS.n2405 5.2005
R3150 VSS.n2400 VSS.n2399 5.2005
R3151 VSS.n2404 VSS.n2400 5.2005
R3152 VSS.n2402 VSS.n2401 5.2005
R3153 VSS.n2403 VSS.n2402 5.2005
R3154 VSS.n412 VSS.n411 5.2005
R3155 VSS.n413 VSS.n412 5.2005
R3156 VSS.n2609 VSS.n2608 5.2005
R3157 VSS.n2608 VSS.n2607 5.2005
R3158 VSS.n2612 VSS.n2611 5.2005
R3159 VSS.n2613 VSS.n2612 5.2005
R3160 VSS.n407 VSS.n406 5.2005
R3161 VSS.n2614 VSS.n407 5.2005
R3162 VSS.n2617 VSS.n2616 5.2005
R3163 VSS.n2616 VSS.n2615 5.2005
R3164 VSS.n2618 VSS.n405 5.2005
R3165 VSS.n405 VSS.n404 5.2005
R3166 VSS.n2620 VSS.n2619 5.2005
R3167 VSS.n2621 VSS.n2620 5.2005
R3168 VSS.n403 VSS.n402 5.2005
R3169 VSS.n2622 VSS.n403 5.2005
R3170 VSS.n2625 VSS.n2624 5.2005
R3171 VSS.n2624 VSS.n2623 5.2005
R3172 VSS.n2626 VSS.n401 5.2005
R3173 VSS.n401 VSS.n400 5.2005
R3174 VSS.n2630 VSS.n2629 5.2005
R3175 VSS.n2631 VSS.n2630 5.2005
R3176 VSS.n399 VSS.n398 5.2005
R3177 VSS.n2632 VSS.n399 5.2005
R3178 VSS.n2635 VSS.n2634 5.2005
R3179 VSS.n2634 VSS.n2633 5.2005
R3180 VSS.n2636 VSS.n397 5.2005
R3181 VSS.n397 VSS.n396 5.2005
R3182 VSS.n2638 VSS.n2637 5.2005
R3183 VSS.n2639 VSS.n2638 5.2005
R3184 VSS.n395 VSS.n394 5.2005
R3185 VSS.n2640 VSS.n395 5.2005
R3186 VSS.n2643 VSS.n2642 5.2005
R3187 VSS.n2642 VSS.n2641 5.2005
R3188 VSS.n2644 VSS.n393 5.2005
R3189 VSS.n393 VSS.n392 5.2005
R3190 VSS.n2646 VSS.n2645 5.2005
R3191 VSS.n2647 VSS.n2646 5.2005
R3192 VSS.n391 VSS.n390 5.2005
R3193 VSS.n2648 VSS.n391 5.2005
R3194 VSS.n2651 VSS.n2650 5.2005
R3195 VSS.n2650 VSS.n2649 5.2005
R3196 VSS.n2707 VSS.n2706 5.2005
R3197 VSS.n2708 VSS.n2707 5.2005
R3198 VSS.n2705 VSS.n381 5.2005
R3199 VSS.n381 VSS.n379 5.2005
R3200 VSS.n2704 VSS.n2703 5.2005
R3201 VSS.n2703 VSS.n2702 5.2005
R3202 VSS.n2654 VSS.n2653 5.2005
R3203 VSS.n2701 VSS.n2654 5.2005
R3204 VSS.n2699 VSS.n2698 5.2005
R3205 VSS.n2700 VSS.n2699 5.2005
R3206 VSS.n2697 VSS.n2656 5.2005
R3207 VSS.n2656 VSS.n2655 5.2005
R3208 VSS.n2696 VSS.n2695 5.2005
R3209 VSS.n2695 VSS.n2694 5.2005
R3210 VSS.n2658 VSS.n2657 5.2005
R3211 VSS.n2693 VSS.n2658 5.2005
R3212 VSS.n2691 VSS.n2690 5.2005
R3213 VSS.n2692 VSS.n2691 5.2005
R3214 VSS.n2688 VSS.n2660 5.2005
R3215 VSS.n2660 VSS.n2659 5.2005
R3216 VSS.n2687 VSS.n2686 5.2005
R3217 VSS.n2686 VSS.n2685 5.2005
R3218 VSS.n2663 VSS.n2662 5.2005
R3219 VSS.n2684 VSS.n2663 5.2005
R3220 VSS.n2682 VSS.n2681 5.2005
R3221 VSS.n2683 VSS.n2682 5.2005
R3222 VSS.n2680 VSS.n2665 5.2005
R3223 VSS.n2665 VSS.n2664 5.2005
R3224 VSS.n2679 VSS.n2678 5.2005
R3225 VSS.n2678 VSS.n2677 5.2005
R3226 VSS.n2667 VSS.n2666 5.2005
R3227 VSS.n2676 VSS.n2667 5.2005
R3228 VSS.n2674 VSS.n2673 5.2005
R3229 VSS.n2675 VSS.n2674 5.2005
R3230 VSS.n2672 VSS.n2669 5.2005
R3231 VSS.n2669 VSS.n2668 5.2005
R3232 VSS.n2671 VSS.n2670 5.2005
R3233 VSS.n2670 VSS.n267 5.2005
R3234 VSS.n2883 VSS.n2882 5.2005
R3235 VSS.n2882 VSS.n2881 5.2005
R3236 VSS.n2884 VSS.n263 5.2005
R3237 VSS.n263 VSS.n262 5.2005
R3238 VSS.n2886 VSS.n2885 5.2005
R3239 VSS.n2887 VSS.n2886 5.2005
R3240 VSS.n261 VSS.n260 5.2005
R3241 VSS.n2888 VSS.n261 5.2005
R3242 VSS.n2891 VSS.n2890 5.2005
R3243 VSS.n2890 VSS.n2889 5.2005
R3244 VSS.n2892 VSS.n259 5.2005
R3245 VSS.n259 VSS.n258 5.2005
R3246 VSS.n2894 VSS.n2893 5.2005
R3247 VSS.n2895 VSS.n2894 5.2005
R3248 VSS.n257 VSS.n256 5.2005
R3249 VSS.n2896 VSS.n257 5.2005
R3250 VSS.n2899 VSS.n2898 5.2005
R3251 VSS.n2898 VSS.n2897 5.2005
R3252 VSS.n2901 VSS.n254 5.2005
R3253 VSS.n254 VSS.n253 5.2005
R3254 VSS.n2903 VSS.n2902 5.2005
R3255 VSS.n2904 VSS.n2903 5.2005
R3256 VSS.n252 VSS.n251 5.2005
R3257 VSS.n2905 VSS.n252 5.2005
R3258 VSS.n2908 VSS.n2907 5.2005
R3259 VSS.n2907 VSS.n2906 5.2005
R3260 VSS.n2909 VSS.n250 5.2005
R3261 VSS.n250 VSS.n249 5.2005
R3262 VSS.n2911 VSS.n2910 5.2005
R3263 VSS.n2912 VSS.n2911 5.2005
R3264 VSS.n248 VSS.n247 5.2005
R3265 VSS.n2913 VSS.n248 5.2005
R3266 VSS.n2916 VSS.n2915 5.2005
R3267 VSS.n2915 VSS.n2914 5.2005
R3268 VSS.n2917 VSS.n245 5.2005
R3269 VSS.n245 VSS.n243 5.2005
R3270 VSS.n2942 VSS.n2941 5.2005
R3271 VSS.n2943 VSS.n2942 5.2005
R3272 VSS.n2939 VSS.n2938 5.2005
R3273 VSS.n2938 VSS.n2937 5.2005
R3274 VSS.n2927 VSS.n2926 5.2005
R3275 VSS.n2936 VSS.n2927 5.2005
R3276 VSS.n2934 VSS.n2933 5.2005
R3277 VSS.n2935 VSS.n2934 5.2005
R3278 VSS.n2932 VSS.n2929 5.2005
R3279 VSS.n2929 VSS.n2928 5.2005
R3280 VSS.n2931 VSS.n2930 5.2005
R3281 VSS.n2930 VSS.n201 5.2005
R3282 VSS.n200 VSS.n199 5.2005
R3283 VSS.n2962 VSS.n200 5.2005
R3284 VSS.n2965 VSS.n2964 5.2005
R3285 VSS.n2964 VSS.n2963 5.2005
R3286 VSS.n2966 VSS.n198 5.2005
R3287 VSS.n198 VSS.n197 5.2005
R3288 VSS.n2969 VSS.n2968 5.2005
R3289 VSS.n2970 VSS.n2969 5.2005
R3290 VSS.n2967 VSS.n196 5.2005
R3291 VSS.n2971 VSS.n196 5.2005
R3292 VSS.n2974 VSS.n2973 5.2005
R3293 VSS.n2973 VSS.n2972 5.2005
R3294 VSS.n2975 VSS.n193 5.2005
R3295 VSS.n193 VSS.n192 5.2005
R3296 VSS.n2977 VSS.n2976 5.2005
R3297 VSS.n2978 VSS.n2977 5.2005
R3298 VSS.n191 VSS.n190 5.2005
R3299 VSS.n2979 VSS.n191 5.2005
R3300 VSS.n2982 VSS.n2981 5.2005
R3301 VSS.n2981 VSS.n2980 5.2005
R3302 VSS.n2983 VSS.n189 5.2005
R3303 VSS.n189 VSS.n188 5.2005
R3304 VSS.n2985 VSS.n2984 5.2005
R3305 VSS.n2986 VSS.n2985 5.2005
R3306 VSS.n187 VSS.n186 5.2005
R3307 VSS.n2987 VSS.n187 5.2005
R3308 VSS.n2990 VSS.n2989 5.2005
R3309 VSS.n2989 VSS.n2988 5.2005
R3310 VSS.n3039 VSS.n3038 5.2005
R3311 VSS.n3040 VSS.n3039 5.2005
R3312 VSS.n3037 VSS.n173 5.2005
R3313 VSS.n173 VSS.n171 5.2005
R3314 VSS.n3036 VSS.n3035 5.2005
R3315 VSS.n3035 VSS.n3034 5.2005
R3316 VSS.n2993 VSS.n2992 5.2005
R3317 VSS.n3033 VSS.n2993 5.2005
R3318 VSS.n3031 VSS.n3030 5.2005
R3319 VSS.n3032 VSS.n3031 5.2005
R3320 VSS.n3029 VSS.n2994 5.2005
R3321 VSS.n3028 VSS.n3027 5.2005
R3322 VSS.n3027 VSS.n3026 5.2005
R3323 VSS.n2996 VSS.n2995 5.2005
R3324 VSS.n3025 VSS.n2996 5.2005
R3325 VSS.n3023 VSS.n3022 5.2005
R3326 VSS.n3024 VSS.n3023 5.2005
R3327 VSS.n3021 VSS.n2999 5.2005
R3328 VSS.n2999 VSS.n2998 5.2005
R3329 VSS.n3020 VSS.n3019 5.2005
R3330 VSS.n3019 VSS.n3018 5.2005
R3331 VSS.n3001 VSS.n3000 5.2005
R3332 VSS.n3017 VSS.n3001 5.2005
R3333 VSS.n3015 VSS.n3014 5.2005
R3334 VSS.n3016 VSS.n3015 5.2005
R3335 VSS.n3013 VSS.n3003 5.2005
R3336 VSS.n3003 VSS.n3002 5.2005
R3337 VSS.n3012 VSS.n3011 5.2005
R3338 VSS.n3011 VSS.n3010 5.2005
R3339 VSS.n3005 VSS.n3004 5.2005
R3340 VSS.n3009 VSS.n3005 5.2005
R3341 VSS.n3007 VSS.n3006 5.2005
R3342 VSS.n3008 VSS.n3007 5.2005
R3343 VSS.n3 VSS.n2 5.2005
R3344 VSS.n5 VSS.n3 5.2005
R3345 VSS.n3483 VSS.n3482 5.2005
R3346 VSS.n3482 VSS.n3481 5.2005
R3347 VSS.n3484 VSS.n3483 5.15774
R3348 VSS VSS.n3484 5.05708
R3349 VSS.n1608 VSS.n1106 4.83445
R3350 VSS.n223 VSS.n119 4.74734
R3351 VSS.n165 VSS.n163 4.51084
R3352 VSS.n3429 VSS.n70 4.50813
R3353 VSS.n1753 VSS.n1007 4.5005
R3354 VSS.n1753 VSS.n1008 4.5005
R3355 VSS.n1753 VSS.n1006 4.5005
R3356 VSS.n1753 VSS.n1009 4.5005
R3357 VSS.n1753 VSS.n1005 4.5005
R3358 VSS.n1753 VSS.n1010 4.5005
R3359 VSS.n1753 VSS.n1004 4.5005
R3360 VSS.n1753 VSS.n1752 4.5005
R3361 VSS.n1024 VSS.n1006 4.5005
R3362 VSS.n1024 VSS.n1009 4.5005
R3363 VSS.n1024 VSS.n1005 4.5005
R3364 VSS.n1024 VSS.n1010 4.5005
R3365 VSS.n1024 VSS.n1004 4.5005
R3366 VSS.n1752 VSS.n1024 4.5005
R3367 VSS.n1024 VSS.n1003 4.5005
R3368 VSS.n1019 VSS.n1006 4.5005
R3369 VSS.n1019 VSS.n1009 4.5005
R3370 VSS.n1019 VSS.n1005 4.5005
R3371 VSS.n1019 VSS.n1010 4.5005
R3372 VSS.n1019 VSS.n1004 4.5005
R3373 VSS.n1752 VSS.n1019 4.5005
R3374 VSS.n1019 VSS.n1003 4.5005
R3375 VSS.n1027 VSS.n1006 4.5005
R3376 VSS.n1027 VSS.n1009 4.5005
R3377 VSS.n1027 VSS.n1005 4.5005
R3378 VSS.n1027 VSS.n1010 4.5005
R3379 VSS.n1027 VSS.n1004 4.5005
R3380 VSS.n1752 VSS.n1027 4.5005
R3381 VSS.n1027 VSS.n1003 4.5005
R3382 VSS.n1018 VSS.n1006 4.5005
R3383 VSS.n1018 VSS.n1009 4.5005
R3384 VSS.n1018 VSS.n1005 4.5005
R3385 VSS.n1018 VSS.n1010 4.5005
R3386 VSS.n1018 VSS.n1004 4.5005
R3387 VSS.n1752 VSS.n1018 4.5005
R3388 VSS.n1018 VSS.n1003 4.5005
R3389 VSS.n1030 VSS.n1006 4.5005
R3390 VSS.n1030 VSS.n1009 4.5005
R3391 VSS.n1030 VSS.n1005 4.5005
R3392 VSS.n1030 VSS.n1010 4.5005
R3393 VSS.n1030 VSS.n1004 4.5005
R3394 VSS.n1752 VSS.n1030 4.5005
R3395 VSS.n1030 VSS.n1003 4.5005
R3396 VSS.n1017 VSS.n1006 4.5005
R3397 VSS.n1017 VSS.n1009 4.5005
R3398 VSS.n1017 VSS.n1005 4.5005
R3399 VSS.n1017 VSS.n1010 4.5005
R3400 VSS.n1017 VSS.n1004 4.5005
R3401 VSS.n1752 VSS.n1017 4.5005
R3402 VSS.n1017 VSS.n1003 4.5005
R3403 VSS.n1033 VSS.n1006 4.5005
R3404 VSS.n1033 VSS.n1009 4.5005
R3405 VSS.n1033 VSS.n1005 4.5005
R3406 VSS.n1033 VSS.n1010 4.5005
R3407 VSS.n1033 VSS.n1004 4.5005
R3408 VSS.n1752 VSS.n1033 4.5005
R3409 VSS.n1033 VSS.n1003 4.5005
R3410 VSS.n1016 VSS.n1006 4.5005
R3411 VSS.n1016 VSS.n1009 4.5005
R3412 VSS.n1016 VSS.n1005 4.5005
R3413 VSS.n1016 VSS.n1010 4.5005
R3414 VSS.n1016 VSS.n1004 4.5005
R3415 VSS.n1752 VSS.n1016 4.5005
R3416 VSS.n1016 VSS.n1003 4.5005
R3417 VSS.n1036 VSS.n1006 4.5005
R3418 VSS.n1036 VSS.n1009 4.5005
R3419 VSS.n1036 VSS.n1005 4.5005
R3420 VSS.n1036 VSS.n1010 4.5005
R3421 VSS.n1036 VSS.n1004 4.5005
R3422 VSS.n1752 VSS.n1036 4.5005
R3423 VSS.n1036 VSS.n1003 4.5005
R3424 VSS.n1015 VSS.n1006 4.5005
R3425 VSS.n1015 VSS.n1009 4.5005
R3426 VSS.n1015 VSS.n1005 4.5005
R3427 VSS.n1015 VSS.n1010 4.5005
R3428 VSS.n1015 VSS.n1004 4.5005
R3429 VSS.n1752 VSS.n1015 4.5005
R3430 VSS.n1015 VSS.n1003 4.5005
R3431 VSS.n1039 VSS.n1006 4.5005
R3432 VSS.n1039 VSS.n1009 4.5005
R3433 VSS.n1039 VSS.n1005 4.5005
R3434 VSS.n1039 VSS.n1010 4.5005
R3435 VSS.n1039 VSS.n1004 4.5005
R3436 VSS.n1752 VSS.n1039 4.5005
R3437 VSS.n1039 VSS.n1003 4.5005
R3438 VSS.n1014 VSS.n1006 4.5005
R3439 VSS.n1014 VSS.n1009 4.5005
R3440 VSS.n1014 VSS.n1005 4.5005
R3441 VSS.n1014 VSS.n1010 4.5005
R3442 VSS.n1014 VSS.n1004 4.5005
R3443 VSS.n1752 VSS.n1014 4.5005
R3444 VSS.n1014 VSS.n1003 4.5005
R3445 VSS.n1042 VSS.n1006 4.5005
R3446 VSS.n1042 VSS.n1009 4.5005
R3447 VSS.n1042 VSS.n1005 4.5005
R3448 VSS.n1042 VSS.n1010 4.5005
R3449 VSS.n1042 VSS.n1004 4.5005
R3450 VSS.n1752 VSS.n1042 4.5005
R3451 VSS.n1042 VSS.n1003 4.5005
R3452 VSS.n1013 VSS.n1006 4.5005
R3453 VSS.n1013 VSS.n1009 4.5005
R3454 VSS.n1013 VSS.n1005 4.5005
R3455 VSS.n1013 VSS.n1010 4.5005
R3456 VSS.n1013 VSS.n1004 4.5005
R3457 VSS.n1752 VSS.n1013 4.5005
R3458 VSS.n1013 VSS.n1003 4.5005
R3459 VSS.n1044 VSS.n1006 4.5005
R3460 VSS.n1044 VSS.n1009 4.5005
R3461 VSS.n1044 VSS.n1005 4.5005
R3462 VSS.n1044 VSS.n1010 4.5005
R3463 VSS.n1044 VSS.n1004 4.5005
R3464 VSS.n1752 VSS.n1044 4.5005
R3465 VSS.n1044 VSS.n1003 4.5005
R3466 VSS.n1045 VSS.n1007 4.5005
R3467 VSS.n1045 VSS.n1008 4.5005
R3468 VSS.n1045 VSS.n1006 4.5005
R3469 VSS.n1045 VSS.n1009 4.5005
R3470 VSS.n1045 VSS.n1005 4.5005
R3471 VSS.n1045 VSS.n1010 4.5005
R3472 VSS.n1045 VSS.n1004 4.5005
R3473 VSS.n1752 VSS.n1045 4.5005
R3474 VSS.n1751 VSS.n1007 4.5005
R3475 VSS.n1751 VSS.n1008 4.5005
R3476 VSS.n1751 VSS.n1006 4.5005
R3477 VSS.n1751 VSS.n1009 4.5005
R3478 VSS.n1751 VSS.n1005 4.5005
R3479 VSS.n1751 VSS.n1010 4.5005
R3480 VSS.n1751 VSS.n1004 4.5005
R3481 VSS.n1752 VSS.n1751 4.5005
R3482 VSS.n1751 VSS.n1003 4.5005
R3483 VSS.n1021 VSS.n1006 4.5005
R3484 VSS.n1021 VSS.n1009 4.5005
R3485 VSS.n1021 VSS.n1005 4.5005
R3486 VSS.n1021 VSS.n1010 4.5005
R3487 VSS.n1021 VSS.n1004 4.5005
R3488 VSS.n1752 VSS.n1021 4.5005
R3489 VSS.n1021 VSS.n1003 4.5005
R3490 VSS.n1008 VSS.n627 4.5005
R3491 VSS.n1006 VSS.n627 4.5005
R3492 VSS.n1009 VSS.n627 4.5005
R3493 VSS.n1005 VSS.n627 4.5005
R3494 VSS.n1010 VSS.n627 4.5005
R3495 VSS.n1004 VSS.n627 4.5005
R3496 VSS.n1752 VSS.n627 4.5005
R3497 VSS.n1003 VSS.n627 4.5005
R3498 VSS.n1753 VSS.n1003 4.5005
R3499 VSS.n1000 VSS.n620 4.5005
R3500 VSS.n999 VSS.n642 4.5005
R3501 VSS.n646 VSS.n641 4.5005
R3502 VSS.n995 VSS.n994 4.5005
R3503 VSS.n993 VSS.n645 4.5005
R3504 VSS.n992 VSS.n991 4.5005
R3505 VSS.n649 VSS.n647 4.5005
R3506 VSS.n987 VSS.n986 4.5005
R3507 VSS.n985 VSS.n652 4.5005
R3508 VSS.n984 VSS.n983 4.5005
R3509 VSS.n667 VSS.n653 4.5005
R3510 VSS.n979 VSS.n978 4.5005
R3511 VSS.n977 VSS.n670 4.5005
R3512 VSS.n976 VSS.n975 4.5005
R3513 VSS.n673 VSS.n671 4.5005
R3514 VSS.n971 VSS.n970 4.5005
R3515 VSS.n969 VSS.n676 4.5005
R3516 VSS.n968 VSS.n967 4.5005
R3517 VSS.n965 VSS.n949 4.5005
R3518 VSS.n1754 VSS.n630 4.5005
R3519 VSS.n1754 VSS.n621 4.5005
R3520 VSS.n1757 VSS.n622 4.5005
R3521 VSS.n1755 VSS.n622 4.5005
R3522 VSS.n1756 VSS.n630 4.5005
R3523 VSS.n1756 VSS.n626 4.5005
R3524 VSS.n1756 VSS.n632 4.5005
R3525 VSS.n1756 VSS.n625 4.5005
R3526 VSS.n1756 VSS.n634 4.5005
R3527 VSS.n1756 VSS.n621 4.5005
R3528 VSS.n1757 VSS.n1756 4.5005
R3529 VSS.n1756 VSS.n1755 4.5005
R3530 VSS.n1755 VSS.n1754 4.5005
R3531 VSS.n1747 VSS.n1721 4.5005
R3532 VSS.n1749 VSS.n1721 4.5005
R3533 VSS.n1717 VSS.n1697 4.5005
R3534 VSS.n1747 VSS.n1717 4.5005
R3535 VSS.n1749 VSS.n1717 4.5005
R3536 VSS.n1723 VSS.n1697 4.5005
R3537 VSS.n1723 VSS.n1053 4.5005
R3538 VSS.n1723 VSS.n1698 4.5005
R3539 VSS.n1723 VSS.n1052 4.5005
R3540 VSS.n1723 VSS.n1699 4.5005
R3541 VSS.n1747 VSS.n1723 4.5005
R3542 VSS.n1749 VSS.n1723 4.5005
R3543 VSS.n1714 VSS.n1697 4.5005
R3544 VSS.n1714 VSS.n1053 4.5005
R3545 VSS.n1714 VSS.n1698 4.5005
R3546 VSS.n1714 VSS.n1052 4.5005
R3547 VSS.n1714 VSS.n1699 4.5005
R3548 VSS.n1747 VSS.n1714 4.5005
R3549 VSS.n1749 VSS.n1714 4.5005
R3550 VSS.n1725 VSS.n1697 4.5005
R3551 VSS.n1725 VSS.n1053 4.5005
R3552 VSS.n1725 VSS.n1698 4.5005
R3553 VSS.n1725 VSS.n1052 4.5005
R3554 VSS.n1725 VSS.n1699 4.5005
R3555 VSS.n1747 VSS.n1725 4.5005
R3556 VSS.n1749 VSS.n1725 4.5005
R3557 VSS.n1713 VSS.n1697 4.5005
R3558 VSS.n1713 VSS.n1053 4.5005
R3559 VSS.n1713 VSS.n1698 4.5005
R3560 VSS.n1713 VSS.n1052 4.5005
R3561 VSS.n1713 VSS.n1699 4.5005
R3562 VSS.n1747 VSS.n1713 4.5005
R3563 VSS.n1749 VSS.n1713 4.5005
R3564 VSS.n1727 VSS.n1697 4.5005
R3565 VSS.n1727 VSS.n1053 4.5005
R3566 VSS.n1727 VSS.n1698 4.5005
R3567 VSS.n1727 VSS.n1052 4.5005
R3568 VSS.n1727 VSS.n1699 4.5005
R3569 VSS.n1747 VSS.n1727 4.5005
R3570 VSS.n1749 VSS.n1727 4.5005
R3571 VSS.n1712 VSS.n1697 4.5005
R3572 VSS.n1712 VSS.n1053 4.5005
R3573 VSS.n1712 VSS.n1698 4.5005
R3574 VSS.n1712 VSS.n1052 4.5005
R3575 VSS.n1712 VSS.n1699 4.5005
R3576 VSS.n1747 VSS.n1712 4.5005
R3577 VSS.n1749 VSS.n1712 4.5005
R3578 VSS.n1729 VSS.n1697 4.5005
R3579 VSS.n1729 VSS.n1053 4.5005
R3580 VSS.n1729 VSS.n1698 4.5005
R3581 VSS.n1729 VSS.n1052 4.5005
R3582 VSS.n1729 VSS.n1699 4.5005
R3583 VSS.n1747 VSS.n1729 4.5005
R3584 VSS.n1749 VSS.n1729 4.5005
R3585 VSS.n1711 VSS.n1697 4.5005
R3586 VSS.n1711 VSS.n1053 4.5005
R3587 VSS.n1711 VSS.n1698 4.5005
R3588 VSS.n1711 VSS.n1052 4.5005
R3589 VSS.n1711 VSS.n1699 4.5005
R3590 VSS.n1747 VSS.n1711 4.5005
R3591 VSS.n1749 VSS.n1711 4.5005
R3592 VSS.n1731 VSS.n1697 4.5005
R3593 VSS.n1731 VSS.n1053 4.5005
R3594 VSS.n1731 VSS.n1698 4.5005
R3595 VSS.n1731 VSS.n1052 4.5005
R3596 VSS.n1731 VSS.n1699 4.5005
R3597 VSS.n1747 VSS.n1731 4.5005
R3598 VSS.n1749 VSS.n1731 4.5005
R3599 VSS.n1710 VSS.n1697 4.5005
R3600 VSS.n1710 VSS.n1053 4.5005
R3601 VSS.n1710 VSS.n1698 4.5005
R3602 VSS.n1710 VSS.n1052 4.5005
R3603 VSS.n1710 VSS.n1699 4.5005
R3604 VSS.n1747 VSS.n1710 4.5005
R3605 VSS.n1749 VSS.n1710 4.5005
R3606 VSS.n1733 VSS.n1697 4.5005
R3607 VSS.n1733 VSS.n1053 4.5005
R3608 VSS.n1733 VSS.n1698 4.5005
R3609 VSS.n1733 VSS.n1052 4.5005
R3610 VSS.n1733 VSS.n1699 4.5005
R3611 VSS.n1747 VSS.n1733 4.5005
R3612 VSS.n1749 VSS.n1733 4.5005
R3613 VSS.n1709 VSS.n1697 4.5005
R3614 VSS.n1709 VSS.n1053 4.5005
R3615 VSS.n1709 VSS.n1698 4.5005
R3616 VSS.n1709 VSS.n1052 4.5005
R3617 VSS.n1709 VSS.n1699 4.5005
R3618 VSS.n1747 VSS.n1709 4.5005
R3619 VSS.n1749 VSS.n1709 4.5005
R3620 VSS.n1735 VSS.n1697 4.5005
R3621 VSS.n1735 VSS.n1053 4.5005
R3622 VSS.n1735 VSS.n1698 4.5005
R3623 VSS.n1735 VSS.n1052 4.5005
R3624 VSS.n1735 VSS.n1699 4.5005
R3625 VSS.n1747 VSS.n1735 4.5005
R3626 VSS.n1749 VSS.n1735 4.5005
R3627 VSS.n1708 VSS.n1697 4.5005
R3628 VSS.n1708 VSS.n1053 4.5005
R3629 VSS.n1708 VSS.n1698 4.5005
R3630 VSS.n1708 VSS.n1052 4.5005
R3631 VSS.n1708 VSS.n1699 4.5005
R3632 VSS.n1747 VSS.n1708 4.5005
R3633 VSS.n1749 VSS.n1708 4.5005
R3634 VSS.n1748 VSS.n1697 4.5005
R3635 VSS.n1748 VSS.n1053 4.5005
R3636 VSS.n1748 VSS.n1698 4.5005
R3637 VSS.n1748 VSS.n1052 4.5005
R3638 VSS.n1748 VSS.n1699 4.5005
R3639 VSS.n1748 VSS.n1747 4.5005
R3640 VSS.n1749 VSS.n1748 4.5005
R3641 VSS.n1702 VSS.n1697 4.5005
R3642 VSS.n1702 VSS.n1053 4.5005
R3643 VSS.n1702 VSS.n1698 4.5005
R3644 VSS.n1702 VSS.n1052 4.5005
R3645 VSS.n1702 VSS.n1699 4.5005
R3646 VSS.n1747 VSS.n1702 4.5005
R3647 VSS.n1749 VSS.n1702 4.5005
R3648 VSS.n1750 VSS.n1697 4.5005
R3649 VSS.n1750 VSS.n1053 4.5005
R3650 VSS.n1750 VSS.n1698 4.5005
R3651 VSS.n1750 VSS.n1052 4.5005
R3652 VSS.n1750 VSS.n1699 4.5005
R3653 VSS.n1750 VSS.n1749 4.5005
R3654 VSS.n3470 VSS.n14 4.43655
R3655 VSS.n2176 VSS.n2175 4.43088
R3656 VSS.n2180 VSS.n2179 4.43088
R3657 VSS.n2181 VSS.n2180 4.43088
R3658 VSS.n2185 VSS.n2184 4.43088
R3659 VSS.n2207 VSS.n2206 4.43088
R3660 VSS.n2204 VSS.n2188 4.43088
R3661 VSS.n2200 VSS.n2199 4.43088
R3662 VSS.n2197 VSS.n2191 4.43088
R3663 VSS.n1471 VSS.n1470 4.43088
R3664 VSS.n1471 VSS.n1462 4.43088
R3665 VSS.n1475 VSS.n1462 4.43088
R3666 VSS.n1475 VSS.n1460 4.43088
R3667 VSS.n1480 VSS.n1460 4.43088
R3668 VSS.n1480 VSS.n1458 4.43088
R3669 VSS.n1484 VSS.n1458 4.43088
R3670 VSS.n1485 VSS.n1484 4.43088
R3671 VSS.n1485 VSS.n1457 4.43088
R3672 VSS.n1489 VSS.n1457 4.43088
R3673 VSS.n1489 VSS.n1455 4.43088
R3674 VSS.n1493 VSS.n1455 4.43088
R3675 VSS.n1493 VSS.n1452 4.43088
R3676 VSS.n1504 VSS.n1452 4.43088
R3677 VSS.n1504 VSS.n1453 4.43088
R3678 VSS.n1500 VSS.n1499 4.43088
R3679 VSS.n165 VSS.n164 4.38259
R3680 VSS.n1393 VSS.n1149 4.33234
R3681 VSS.t100 VSS.t104 4.27307
R3682 VSS.n1362 VSS.n1218 4.13154
R3683 VSS.n1660 VSS.n1063 4.12546
R3684 VSS.n1663 VSS.n1063 4.12546
R3685 VSS.n3446 VSS.n26 4.11885
R3686 VSS.n1573 VSS.t37 4.0955
R3687 VSS.n1572 VSS.t161 4.0955
R3688 VSS.n1420 VSS.t172 4.0955
R3689 VSS.n2304 VSS.n2303 4.05793
R3690 VSS.n2463 VSS.n476 4.05793
R3691 VSS.n2571 VSS.n2570 4.05793
R3692 VSS.n2746 VSS.n354 4.05793
R3693 VSS.n2843 VSS.n2842 4.05793
R3694 VSS.n1409 VSS.t202 4.04494
R3695 VSS.n1409 VSS.t206 4.04494
R3696 VSS.n1577 VSS.t197 4.04494
R3697 VSS.n1577 VSS.t208 4.04494
R3698 VSS.n1576 VSS.t107 4.04494
R3699 VSS.n1576 VSS.t209 4.04494
R3700 VSS.n1417 VSS.t20 4.04494
R3701 VSS.n1417 VSS.t204 4.04494
R3702 VSS.n1590 VSS.n1415 3.89923
R3703 VSS.n1079 VSS.n597 3.8975
R3704 VSS.n1560 VSS.t244 3.8098
R3705 VSS.n1560 VSS.t248 3.8098
R3706 VSS.n1561 VSS.t236 3.8098
R3707 VSS.n1561 VSS.t246 3.8098
R3708 VSS.n1562 VSS.t250 3.8098
R3709 VSS.n1562 VSS.t238 3.8098
R3710 VSS.n1689 VSS.n1688 3.80605
R3711 VSS.n1684 VSS.n1069 3.80605
R3712 VSS.n1680 VSS.n1068 3.80605
R3713 VSS.n1676 VSS.n1067 3.80605
R3714 VSS.n1672 VSS.n1066 3.80605
R3715 VSS.n1668 VSS.n1065 3.80605
R3716 VSS.n1664 VSS.n1064 3.80605
R3717 VSS.n1667 VSS.n1064 3.80605
R3718 VSS.n1671 VSS.n1065 3.80605
R3719 VSS.n1675 VSS.n1066 3.80605
R3720 VSS.n1679 VSS.n1067 3.80605
R3721 VSS.n1683 VSS.n1068 3.80605
R3722 VSS.n1070 VSS.n1069 3.80605
R3723 VSS.n1689 VSS.n1060 3.80605
R3724 VSS.n1200 VSS.n1163 3.79267
R3725 VSS.n1198 VSS.n1166 3.79267
R3726 VSS.n1194 VSS.n1193 3.79267
R3727 VSS.n1187 VSS.n1168 3.79267
R3728 VSS.n1186 VSS.n1185 3.79267
R3729 VSS.n1179 VSS.n1170 3.79267
R3730 VSS.n1178 VSS.n1177 3.79267
R3731 VSS.n1173 VSS.n1172 3.79267
R3732 VSS.n1339 VSS.n1236 3.79267
R3733 VSS.n1335 VSS.n1235 3.79267
R3734 VSS.n1331 VSS.n1234 3.79267
R3735 VSS.n1327 VSS.n1233 3.79267
R3736 VSS.n1323 VSS.n1232 3.79267
R3737 VSS.n1319 VSS.n1231 3.79267
R3738 VSS.n1315 VSS.n1230 3.79267
R3739 VSS.n1311 VSS.n1229 3.79267
R3740 VSS.n1201 VSS.n1200 3.79267
R3741 VSS.n1195 VSS.n1166 3.79267
R3742 VSS.n1193 VSS.n1192 3.79267
R3743 VSS.n1188 VSS.n1187 3.79267
R3744 VSS.n1185 VSS.n1184 3.79267
R3745 VSS.n1180 VSS.n1179 3.79267
R3746 VSS.n1177 VSS.n1176 3.79267
R3747 VSS.n1172 VSS.n1159 3.79267
R3748 VSS.n1314 VSS.n1229 3.79267
R3749 VSS.n1318 VSS.n1230 3.79267
R3750 VSS.n1322 VSS.n1231 3.79267
R3751 VSS.n1326 VSS.n1232 3.79267
R3752 VSS.n1330 VSS.n1233 3.79267
R3753 VSS.n1334 VSS.n1234 3.79267
R3754 VSS.n1338 VSS.n1235 3.79267
R3755 VSS.n1237 VSS.n1236 3.79267
R3756 VSS.n3448 VSS.n3447 3.73488
R3757 VSS.n2302 VSS.n553 3.71266
R3758 VSS.n2091 VSS.n466 3.71266
R3759 VSS.n2569 VSS.n433 3.71266
R3760 VSS.n2747 VSS.n311 3.71266
R3761 VSS.n325 VSS.n99 3.71266
R3762 VSS.t69 VSS.t203 3.71055
R3763 VSS.n3449 VSS.n41 3.69405
R3764 VSS.n3457 VSS.n27 3.69405
R3765 VSS.n3462 VSS.n3461 3.69405
R3766 VSS.n1366 VSS.n1365 3.64321
R3767 VSS.n1365 VSS.n1211 3.64321
R3768 VSS.n1410 VSS.t55 3.6005
R3769 VSS.n1410 VSS.t51 3.6005
R3770 VSS.n291 VSS.n290 3.59261
R3771 VSS.n1921 VSS.n360 3.59261
R3772 VSS.n1862 VSS.n437 3.59261
R3773 VSS.n1782 VSS.n558 3.59261
R3774 VSS.n474 VSS.n467 3.59261
R3775 VSS.n713 VSS.n126 3.59261
R3776 VSS.n812 VSS.n795 3.59261
R3777 VSS.n1097 VSS.t26 3.37782
R3778 VSS.n566 VSS.n565 3.32459
R3779 VSS.n563 VSS.n561 3.32459
R3780 VSS.n2338 VSS.n2337 3.32459
R3781 VSS.n2333 VSS.n535 3.32459
R3782 VSS.n478 VSS.n477 3.32459
R3783 VSS.n2469 VSS.n2468 3.32459
R3784 VSS.n504 VSS.n503 3.32459
R3785 VSS.n507 VSS.n506 3.32459
R3786 VSS.n445 VSS.n444 3.32459
R3787 VSS.n442 VSS.n440 3.32459
R3788 VSS.n2605 VSS.n2604 3.32459
R3789 VSS.n2600 VSS.n415 3.32459
R3790 VSS.n2744 VSS.n2743 3.32459
R3791 VSS.n2739 VSS.n358 3.32459
R3792 VSS.n384 VSS.n377 3.32459
R3793 VSS.n387 VSS.n386 3.32459
R3794 VSS.n2840 VSS.n2839 3.32459
R3795 VSS.n2835 VSS.n288 3.32459
R3796 VSS.n2878 VSS.n2877 3.32459
R3797 VSS.n2873 VSS.n268 3.32459
R3798 VSS.n830 VSS.n829 3.32459
R3799 VSS.n827 VSS.n815 3.32459
R3800 VSS.n823 VSS.n822 3.32459
R3801 VSS.n818 VSS.n817 3.32459
R3802 VSS.n3043 VSS.n3042 3.32459
R3803 VSS.n174 VSS.n170 3.32459
R3804 VSS.n178 VSS.n169 3.32459
R3805 VSS.n182 VSS.n168 3.32459
R3806 VSS.n324 VSS.n321 3.32459
R3807 VSS.n326 VSS.n318 3.32459
R3808 VSS.n348 VSS.n317 3.32459
R3809 VSS.n344 VSS.n316 3.32459
R3810 VSS.n340 VSS.n315 3.32459
R3811 VSS.n336 VSS.n314 3.32459
R3812 VSS.n332 VSS.n286 3.32459
R3813 VSS.n291 VSS.n287 3.32459
R3814 VSS.n1948 VSS.n1913 3.32459
R3815 VSS.n1946 VSS.n1945 3.32459
R3816 VSS.n1940 VSS.n1939 3.32459
R3817 VSS.n1937 VSS.n1936 3.32459
R3818 VSS.n1932 VSS.n1919 3.32459
R3819 VSS.n1930 VSS.n1929 3.32459
R3820 VSS.n1925 VSS.n356 3.32459
R3821 VSS.n1921 VSS.n357 3.32459
R3822 VSS.n1889 VSS.n1888 3.32459
R3823 VSS.n1886 VSS.n1885 3.32459
R3824 VSS.n1880 VSS.n1879 3.32459
R3825 VSS.n1877 VSS.n1876 3.32459
R3826 VSS.n1872 VSS.n1858 3.32459
R3827 VSS.n1870 VSS.n1869 3.32459
R3828 VSS.n1865 VSS.n1861 3.32459
R3829 VSS.n1863 VSS.n1862 3.32459
R3830 VSS.n1887 VSS.n1886 3.32459
R3831 VSS.n1890 VSS.n1889 3.32459
R3832 VSS.n1947 VSS.n1946 3.32459
R3833 VSS.n1913 VSS.n1910 3.32459
R3834 VSS.n327 VSS.n326 3.32459
R3835 VSS.n324 VSS.n323 3.32459
R3836 VSS.n1808 VSS.n1770 3.32459
R3837 VSS.n1807 VSS.n1806 3.32459
R3838 VSS.n1800 VSS.n1799 3.32459
R3839 VSS.n1797 VSS.n1796 3.32459
R3840 VSS.n1792 VSS.n1778 3.32459
R3841 VSS.n1790 VSS.n1789 3.32459
R3842 VSS.n1785 VSS.n1781 3.32459
R3843 VSS.n1783 VSS.n1782 3.32459
R3844 VSS.n1806 VSS.n1805 3.32459
R3845 VSS.n1809 VSS.n1808 3.32459
R3846 VSS.n1791 VSS.n1790 3.32459
R3847 VSS.n1778 VSS.n1776 3.32459
R3848 VSS.n1798 VSS.n1797 3.32459
R3849 VSS.n1801 VSS.n1800 3.32459
R3850 VSS.n1871 VSS.n1870 3.32459
R3851 VSS.n1858 VSS.n1856 3.32459
R3852 VSS.n1878 VSS.n1877 3.32459
R3853 VSS.n1881 VSS.n1880 3.32459
R3854 VSS.n1931 VSS.n1930 3.32459
R3855 VSS.n1919 VSS.n1917 3.32459
R3856 VSS.n1938 VSS.n1937 3.32459
R3857 VSS.n1941 VSS.n1940 3.32459
R3858 VSS.n339 VSS.n314 3.32459
R3859 VSS.n343 VSS.n315 3.32459
R3860 VSS.n347 VSS.n316 3.32459
R3861 VSS.n319 VSS.n317 3.32459
R3862 VSS.n3042 VSS.n166 3.32459
R3863 VSS.n177 VSS.n170 3.32459
R3864 VSS.n181 VSS.n169 3.32459
R3865 VSS.n184 VSS.n168 3.32459
R3866 VSS.n2878 VSS.n269 3.32459
R3867 VSS.n2871 VSS.n268 3.32459
R3868 VSS.n385 VSS.n384 3.32459
R3869 VSS.n388 VSS.n387 3.32459
R3870 VSS.n2605 VSS.n416 3.32459
R3871 VSS.n415 VSS.n414 3.32459
R3872 VSS.n505 VSS.n504 3.32459
R3873 VSS.n508 VSS.n507 3.32459
R3874 VSS.n2338 VSS.n536 3.32459
R3875 VSS.n535 VSS.n534 3.32459
R3876 VSS.n2840 VSS.n289 3.32459
R3877 VSS.n288 VSS.n284 3.32459
R3878 VSS.n2744 VSS.n359 3.32459
R3879 VSS.n2737 VSS.n358 3.32459
R3880 VSS.n444 VSS.n443 3.32459
R3881 VSS.n440 VSS.n431 3.32459
R3882 VSS.n480 VSS.n478 3.32459
R3883 VSS.n2469 VSS.n479 3.32459
R3884 VSS.n565 VSS.n564 3.32459
R3885 VSS.n561 VSS.n551 3.32459
R3886 VSS.n1784 VSS.n1783 3.32459
R3887 VSS.n1781 VSS.n1779 3.32459
R3888 VSS.n1864 VSS.n1863 3.32459
R3889 VSS.n1861 VSS.n1859 3.32459
R3890 VSS.n1924 VSS.n357 3.32459
R3891 VSS.n1920 VSS.n356 3.32459
R3892 VSS.n331 VSS.n287 3.32459
R3893 VSS.n335 VSS.n286 3.32459
R3894 VSS.n2058 VSS.n2053 3.32459
R3895 VSS.n2090 VSS.n2089 3.32459
R3896 VSS.n2084 VSS.n2083 3.32459
R3897 VSS.n2081 VSS.n2080 3.32459
R3898 VSS.n2076 VSS.n2065 3.32459
R3899 VSS.n2074 VSS.n2073 3.32459
R3900 VSS.n2066 VSS.n473 3.32459
R3901 VSS.n2068 VSS.n475 3.32459
R3902 VSS.n475 VSS.n474 3.32459
R3903 VSS.n2069 VSS.n473 3.32459
R3904 VSS.n2075 VSS.n2074 3.32459
R3905 VSS.n2065 VSS.n2063 3.32459
R3906 VSS.n2082 VSS.n2081 3.32459
R3907 VSS.n2085 VSS.n2084 3.32459
R3908 VSS.n2090 VSS.n2054 3.32459
R3909 VSS.n2056 VSS.n2053 3.32459
R3910 VSS.n757 VSS.n756 3.32459
R3911 VSS.n761 VSS.n760 3.32459
R3912 VSS.n767 VSS.n766 3.32459
R3913 VSS.n773 VSS.n772 3.32459
R3914 VSS.n776 VSS.n775 3.32459
R3915 VSS.n781 VSS.n780 3.32459
R3916 VSS.n909 VSS.n908 3.32459
R3917 VSS.n914 VSS.n913 3.32459
R3918 VSS.n917 VSS.n916 3.32459
R3919 VSS.n922 VSS.n921 3.32459
R3920 VSS.n925 VSS.n924 3.32459
R3921 VSS.n930 VSS.n929 3.32459
R3922 VSS.n933 VSS.n932 3.32459
R3923 VSS.n938 VSS.n937 3.32459
R3924 VSS.n941 VSS.n940 3.32459
R3925 VSS.n740 VSS.n739 3.32459
R3926 VSS.n737 VSS.n736 3.32459
R3927 VSS.n731 VSS.n730 3.32459
R3928 VSS.n728 VSS.n727 3.32459
R3929 VSS.n723 VSS.n709 3.32459
R3930 VSS.n721 VSS.n720 3.32459
R3931 VSS.n716 VSS.n712 3.32459
R3932 VSS.n714 VSS.n713 3.32459
R3933 VSS.n715 VSS.n714 3.32459
R3934 VSS.n712 VSS.n710 3.32459
R3935 VSS.n722 VSS.n721 3.32459
R3936 VSS.n709 VSS.n707 3.32459
R3937 VSS.n729 VSS.n728 3.32459
R3938 VSS.n732 VSS.n731 3.32459
R3939 VSS.n738 VSS.n737 3.32459
R3940 VSS.n741 VSS.n740 3.32459
R3941 VSS.n215 VSS.n214 3.32459
R3942 VSS.n220 VSS.n219 3.32459
R3943 VSS.n2920 VSS.n241 3.32459
R3944 VSS.n2923 VSS.n2922 3.32459
R3945 VSS.n216 VSS.n215 3.32459
R3946 VSS.n221 VSS.n220 3.32459
R3947 VSS.n2921 VSS.n2920 3.32459
R3948 VSS.n2924 VSS.n2923 3.32459
R3949 VSS.n3085 VSS.n3084 3.32459
R3950 VSS.n3082 VSS.n3081 3.32459
R3951 VSS.n858 VSS.n844 3.32459
R3952 VSS.n856 VSS.n855 3.32459
R3953 VSS.n851 VSS.n846 3.32459
R3954 VSS.n895 VSS.n894 3.32459
R3955 VSS.n803 VSS.n802 3.32459
R3956 VSS.n804 VSS.n798 3.32459
R3957 VSS.n811 VSS.n810 3.32459
R3958 VSS.n810 VSS.n809 3.32459
R3959 VSS.n805 VSS.n804 3.32459
R3960 VSS.n802 VSS.n801 3.32459
R3961 VSS.n896 VSS.n895 3.32459
R3962 VSS.n829 VSS.n828 3.32459
R3963 VSS.n824 VSS.n815 3.32459
R3964 VSS.n822 VSS.n821 3.32459
R3965 VSS.n817 VSS.n153 3.32459
R3966 VSS.n846 VSS.n845 3.32459
R3967 VSS.n857 VSS.n856 3.32459
R3968 VSS.n844 VSS.n842 3.32459
R3969 VSS.n3083 VSS.n3082 3.32459
R3970 VSS.n3086 VSS.n3085 3.32459
R3971 VSS.n758 VSS.n757 3.32459
R3972 VSS.n760 VSS.n694 3.32459
R3973 VSS.n768 VSS.n767 3.32459
R3974 VSS.n774 VSS.n773 3.32459
R3975 VSS.n775 VSS.n690 3.32459
R3976 VSS.n782 VSS.n781 3.32459
R3977 VSS.n908 VSS.n687 3.32459
R3978 VSS.n915 VSS.n914 3.32459
R3979 VSS.n916 VSS.n685 3.32459
R3980 VSS.n923 VSS.n922 3.32459
R3981 VSS.n924 VSS.n683 3.32459
R3982 VSS.n931 VSS.n930 3.32459
R3983 VSS.n932 VSS.n681 3.32459
R3984 VSS.n939 VSS.n938 3.32459
R3985 VSS.n940 VSS.n679 3.32459
R3986 VSS.n1610 VSS.n1609 3.25471
R3987 VSS.n3457 VSS.n3456 3.25471
R3988 VSS.n3461 VSS.n23 3.25471
R3989 VSS.n3471 VSS.n3470 3.25471
R3990 VSS.n1567 VSS.n1106 3.22345
R3991 VSS.n1149 VSS.n1148 3.20971
R3992 VSS.n1610 VSS.n1096 3.20971
R3993 VSS.n2216 VSS.n588 3.18236
R3994 VSS.n3443 VSS.n42 3.11113
R3995 VSS.t71 VSS.n1153 3.00489
R3996 VSS.n3473 VSS.n3472 2.91603
R3997 VSS.n1464 VSS.n592 2.72518
R3998 VSS.n1439 VSS.n1438 2.66271
R3999 VSS.n1586 VSS.n1412 2.66171
R4000 VSS.n3450 VSS.n39 2.60721
R4001 VSS.n1250 VSS.n1242 2.54316
R4002 VSS.n1249 VSS.n1247 2.54316
R4003 VSS.n1244 VSS.n1242 2.54316
R4004 VSS.n1633 VSS.t321 2.5205
R4005 VSS.n1633 VSS.t195 2.5205
R4006 VSS.n3465 VSS.n20 2.4855
R4007 VSS.n1690 VSS.n1062 2.38689
R4008 VSS.n1000 VSS.n636 2.2505
R4009 VSS.n999 VSS.n998 2.2505
R4010 VSS.n997 VSS.n641 2.2505
R4011 VSS.n996 VSS.n995 2.2505
R4012 VSS.n645 VSS.n643 2.2505
R4013 VSS.n991 VSS.n990 2.2505
R4014 VSS.n989 VSS.n649 2.2505
R4015 VSS.n988 VSS.n987 2.2505
R4016 VSS.n652 VSS.n650 2.2505
R4017 VSS.n983 VSS.n982 2.2505
R4018 VSS.n981 VSS.n667 2.2505
R4019 VSS.n980 VSS.n979 2.2505
R4020 VSS.n670 VSS.n668 2.2505
R4021 VSS.n975 VSS.n974 2.2505
R4022 VSS.n973 VSS.n673 2.2505
R4023 VSS.n972 VSS.n971 2.2505
R4024 VSS.n676 VSS.n674 2.2505
R4025 VSS.n1707 VSS.n1705 2.25002
R4026 VSS.n1707 VSS.n1704 2.25002
R4027 VSS.n1707 VSS.n1703 2.25002
R4028 VSS.n1707 VSS.n1012 2.25002
R4029 VSS.n1050 VSS.n1047 2.25002
R4030 VSS.n1050 VSS.n1048 2.25002
R4031 VSS.n1050 VSS.n1049 2.25002
R4032 VSS.n1050 VSS.n1011 2.25002
R4033 VSS.n1721 VSS.n1720 2.24986
R4034 VSS.n1721 VSS.n1719 2.24986
R4035 VSS.n1738 VSS.n1721 2.24986
R4036 VSS.n1717 VSS.n1716 2.24986
R4037 VSS.n1717 VSS.n1715 2.24986
R4038 VSS.n1750 VSS.n1700 2.24986
R4039 VSS.n1022 VSS.n1007 2.24873
R4040 VSS.n1026 VSS.n1008 2.24873
R4041 VSS.n1025 VSS.n1007 2.24873
R4042 VSS.n1029 VSS.n1008 2.24873
R4043 VSS.n1028 VSS.n1007 2.24873
R4044 VSS.n1032 VSS.n1008 2.24873
R4045 VSS.n1031 VSS.n1007 2.24873
R4046 VSS.n1035 VSS.n1008 2.24873
R4047 VSS.n1034 VSS.n1007 2.24873
R4048 VSS.n1038 VSS.n1008 2.24873
R4049 VSS.n1037 VSS.n1007 2.24873
R4050 VSS.n1041 VSS.n1008 2.24873
R4051 VSS.n1040 VSS.n1007 2.24873
R4052 VSS.n1043 VSS.n1008 2.24873
R4053 VSS.n1706 VSS.n1007 2.24873
R4054 VSS.n1046 VSS.n1003 2.24873
R4055 VSS.n1020 VSS.n1007 2.24873
R4056 VSS.n1023 VSS.n1008 2.24873
R4057 VSS.n635 VSS.n624 2.24873
R4058 VSS.n1718 VSS.n1701 2.24873
R4059 VSS.n1746 VSS.n1745 2.24873
R4060 VSS.n1722 VSS.n1701 2.24873
R4061 VSS.n1746 VSS.n1744 2.24873
R4062 VSS.n1724 VSS.n1701 2.24873
R4063 VSS.n1746 VSS.n1743 2.24873
R4064 VSS.n1726 VSS.n1701 2.24873
R4065 VSS.n1746 VSS.n1742 2.24873
R4066 VSS.n1728 VSS.n1701 2.24873
R4067 VSS.n1746 VSS.n1741 2.24873
R4068 VSS.n1730 VSS.n1701 2.24873
R4069 VSS.n1746 VSS.n1740 2.24873
R4070 VSS.n1732 VSS.n1701 2.24873
R4071 VSS.n1746 VSS.n1739 2.24873
R4072 VSS.n1734 VSS.n1701 2.24873
R4073 VSS.n1746 VSS.n1737 2.24873
R4074 VSS.n1736 VSS.n1701 2.24873
R4075 VSS.n1746 VSS.n1051 2.24873
R4076 VSS.n1754 VSS.n638 2.24231
R4077 VSS.n1754 VSS.n637 2.24231
R4078 VSS.n1754 VSS.n623 2.24231
R4079 VSS.n629 VSS.n622 2.24231
R4080 VSS.n631 VSS.n622 2.24231
R4081 VSS.n633 VSS.n622 2.24231
R4082 VSS.n948 VSS.n678 2.219
R4083 VSS.n1759 VSS.n619 2.15937
R4084 VSS.n2149 VSS.n613 2.12174
R4085 VSS.n1243 VSS.t3 2.05866
R4086 VSS.n677 VSS.n68 1.99927
R4087 VSS.n1397 VSS.t329 1.99806
R4088 VSS.n1397 VSS.t277 1.99806
R4089 VSS.n1100 VSS.t122 1.99806
R4090 VSS.n1100 VSS.t75 1.99806
R4091 VSS.n1099 VSS.t281 1.99806
R4092 VSS.n1099 VSS.t174 1.99806
R4093 VSS.n1243 VSS.t1 1.96984
R4094 VSS.n1384 VSS.t42 1.87824
R4095 VSS.n1556 VSS.n1445 1.82428
R4096 VSS.n1556 VSS.n1444 1.82428
R4097 VSS.n1469 VSS.n591 1.82428
R4098 VSS.n1463 VSS.n591 1.82428
R4099 VSS.n2192 VSS.n591 1.82428
R4100 VSS.n2198 VSS.n591 1.82428
R4101 VSS.n2190 VSS.n589 1.82428
R4102 VSS.n2205 VSS.n589 1.82428
R4103 VSS.n2186 VSS.n589 1.82428
R4104 VSS.n598 VSS.n589 1.82428
R4105 VSS.n2173 VSS.n600 1.82428
R4106 VSS.n2174 VSS.n2173 1.82428
R4107 VSS.n3044 VSS.n165 1.81881
R4108 VSS.n1413 VSS.n597 1.80163
R4109 VSS.n1055 VSS.n1054 1.7498
R4110 VSS.n2193 VSS.n592 1.7062
R4111 VSS.n1630 VSS.t7 1.6385
R4112 VSS.n1630 VSS.t346 1.6385
R4113 VSS.n1628 VSS.t293 1.6385
R4114 VSS.n1628 VSS.t323 1.6385
R4115 VSS.n1609 VSS.n1608 1.58024
R4116 VSS.n23 VSS.n13 1.58024
R4117 VSS.n3471 VSS.n13 1.58024
R4118 VSS.n3473 VSS.n12 1.58024
R4119 VSS.n2175 VSS.n2174 1.55443
R4120 VSS.n2179 VSS.n600 1.55443
R4121 VSS.n2184 VSS.n598 1.55443
R4122 VSS.n2207 VSS.n2186 1.55443
R4123 VSS.n2205 VSS.n2204 1.55443
R4124 VSS.n2200 VSS.n2190 1.55443
R4125 VSS.n2198 VSS.n2197 1.55443
R4126 VSS.n2193 VSS.n2192 1.55443
R4127 VSS.n1463 VSS.n1415 1.55443
R4128 VSS.n1470 VSS.n1469 1.55443
R4129 VSS.n1500 VSS.n1444 1.55443
R4130 VSS.n1496 VSS.n1445 1.55443
R4131 VSS.n1499 VSS.n1445 1.55443
R4132 VSS.n1453 VSS.n1444 1.55443
R4133 VSS.n1469 VSS.n1416 1.55443
R4134 VSS.n1464 VSS.n1463 1.55443
R4135 VSS.n2192 VSS.n2191 1.55443
R4136 VSS.n2199 VSS.n2198 1.55443
R4137 VSS.n2190 VSS.n2188 1.55443
R4138 VSS.n2206 VSS.n2205 1.55443
R4139 VSS.n2186 VSS.n2185 1.55443
R4140 VSS.n2181 VSS.n598 1.55443
R4141 VSS.n2176 VSS.n600 1.55443
R4142 VSS.n2174 VSS.n602 1.55443
R4143 VSS.n604 VSS.n602 1.55113
R4144 VSS.n1071 VSS.n1055 1.52481
R4145 VSS.n1002 VSS.n1001 1.5005
R4146 VSS.n666 VSS.t338 1.5005
R4147 VSS.n654 VSS.n640 1.5005
R4148 VSS.n656 VSS.n655 1.5005
R4149 VSS.n657 VSS.n644 1.5005
R4150 VSS.n659 VSS.n658 1.5005
R4151 VSS.n660 VSS.n648 1.5005
R4152 VSS.n662 VSS.n661 1.5005
R4153 VSS.n663 VSS.n651 1.5005
R4154 VSS.n665 VSS.n664 1.5005
R4155 VSS.n952 VSS.n951 1.5005
R4156 VSS.n953 VSS.n669 1.5005
R4157 VSS.n955 VSS.n954 1.5005
R4158 VSS.n956 VSS.n672 1.5005
R4159 VSS.n958 VSS.n957 1.5005
R4160 VSS.n959 VSS.n675 1.5005
R4161 VSS.n961 VSS.n960 1.5005
R4162 VSS.n962 VSS.n950 1.5005
R4163 VSS.n964 VSS.n963 1.5005
R4164 VSS.n1001 VSS.n1000 1.5005
R4165 VSS.n999 VSS.n640 1.5005
R4166 VSS.n655 VSS.n641 1.5005
R4167 VSS.n995 VSS.n644 1.5005
R4168 VSS.n658 VSS.n645 1.5005
R4169 VSS.n991 VSS.n648 1.5005
R4170 VSS.n661 VSS.n649 1.5005
R4171 VSS.n987 VSS.n651 1.5005
R4172 VSS.n665 VSS.n652 1.5005
R4173 VSS.n983 VSS.n666 1.5005
R4174 VSS.n951 VSS.n667 1.5005
R4175 VSS.n979 VSS.n669 1.5005
R4176 VSS.n954 VSS.n670 1.5005
R4177 VSS.n975 VSS.n672 1.5005
R4178 VSS.n957 VSS.n673 1.5005
R4179 VSS.n971 VSS.n675 1.5005
R4180 VSS.n960 VSS.n676 1.5005
R4181 VSS.n967 VSS.n950 1.5005
R4182 VSS.n965 VSS.n964 1.5005
R4183 VSS.n3274 VSS.n3273 1.5005
R4184 VSS.n3272 VSS.n3237 1.5005
R4185 VSS.n3271 VSS.n3270 1.5005
R4186 VSS.n3269 VSS.n3238 1.5005
R4187 VSS.n3268 VSS.n3267 1.5005
R4188 VSS.n3266 VSS.n3239 1.5005
R4189 VSS.n3265 VSS.n3264 1.5005
R4190 VSS.n3263 VSS.n3240 1.5005
R4191 VSS.n3262 VSS.n3261 1.5005
R4192 VSS.n3260 VSS.n3241 1.5005
R4193 VSS.n3259 VSS.n3258 1.5005
R4194 VSS.n3257 VSS.n3242 1.5005
R4195 VSS.n3256 VSS.n3255 1.5005
R4196 VSS.n3254 VSS.n3243 1.5005
R4197 VSS.n3253 VSS.n3252 1.5005
R4198 VSS.n3251 VSS.n3244 1.5005
R4199 VSS.n3250 VSS.n3249 1.5005
R4200 VSS.n3248 VSS.n3245 1.5005
R4201 VSS.n3247 VSS.n3246 1.5005
R4202 VSS.n44 VSS.n43 1.5005
R4203 VSS.n2171 VSS.n604 1.45165
R4204 VSS.n1109 VSS.n1089 1.45008
R4205 VSS.t220 VSS.t276 1.41109
R4206 VSS.n1357 VSS.n1356 1.39283
R4207 VSS.n3456 VSS.n28 1.33629
R4208 VSS.n35 VSS.n23 1.33629
R4209 VSS.n35 VSS.n12 1.33629
R4210 VSS.n3472 VSS.n3471 1.33629
R4211 VSS.n946 VSS.n38 1.33022
R4212 VSS.n1247 VSS.n1246 1.32992
R4213 VSS.n1246 VSS.n1242 1.32992
R4214 VSS.n1593 VSS.n1592 1.28295
R4215 VSS.n619 VSS.n618 1.2567
R4216 VSS.n618 VSS.n617 1.25289
R4217 VSS.n2171 VSS.n605 1.18996
R4218 VSS.n2167 VSS.n605 1.18996
R4219 VSS.n2167 VSS.n2166 1.18996
R4220 VSS.n2166 VSS.n607 1.18996
R4221 VSS.n2162 VSS.n607 1.18996
R4222 VSS.n2162 VSS.n609 1.18996
R4223 VSS.n2158 VSS.n609 1.18996
R4224 VSS.n2158 VSS.n612 1.18996
R4225 VSS.n2150 VSS.n1760 1.18996
R4226 VSS.n2146 VSS.n1760 1.18996
R4227 VSS.n2146 VSS.n1763 1.18996
R4228 VSS.n2142 VSS.n1763 1.18996
R4229 VSS.n2142 VSS.n1766 1.18996
R4230 VSS.n2138 VSS.n1766 1.18996
R4231 VSS.n2138 VSS.n1768 1.18996
R4232 VSS.n2134 VSS.n1768 1.18996
R4233 VSS.n2134 VSS.n2131 1.18996
R4234 VSS.n1642 VSS.n1082 1.16769
R4235 VSS.n966 VSS.n674 1.16259
R4236 VSS.n848 VSS.n847 1.16247
R4237 VSS.n3477 VSS.n7 1.16216
R4238 VSS.n66 VSS.n65 1.1255
R4239 VSS.n3407 VSS.n3406 1.1255
R4240 VSS.n3413 VSS.n3408 1.1255
R4241 VSS.n3414 VSS.n63 1.1255
R4242 VSS.n3415 VSS.n64 1.1255
R4243 VSS.n3403 VSS.n3402 1.1255
R4244 VSS.n3422 VSS.n3421 1.1255
R4245 VSS.n3423 VSS.n3170 1.1255
R4246 VSS.n3425 VSS.n3424 1.1255
R4247 VSS.n3401 VSS.n61 1.1255
R4248 VSS.n3400 VSS.n62 1.1255
R4249 VSS.n3177 VSS.n3171 1.1255
R4250 VSS.n3178 VSS.n3175 1.1255
R4251 VSS.n3392 VSS.n3391 1.1255
R4252 VSS.n3390 VSS.n3176 1.1255
R4253 VSS.n3389 VSS.n3388 1.1255
R4254 VSS.n3179 VSS.n59 1.1255
R4255 VSS.n3382 VSS.n60 1.1255
R4256 VSS.n3381 VSS.n3380 1.1255
R4257 VSS.n3379 VSS.n3183 1.1255
R4258 VSS.n3378 VSS.n3377 1.1255
R4259 VSS.n3185 VSS.n3184 1.1255
R4260 VSS.n3188 VSS.n57 1.1255
R4261 VSS.n3191 VSS.n58 1.1255
R4262 VSS.n3366 VSS.n3365 1.1255
R4263 VSS.n3364 VSS.n3192 1.1255
R4264 VSS.n3363 VSS.n3362 1.1255
R4265 VSS.n3194 VSS.n3193 1.1255
R4266 VSS.n3356 VSS.n3355 1.1255
R4267 VSS.n3354 VSS.n55 1.1255
R4268 VSS.n3353 VSS.n56 1.1255
R4269 VSS.n3202 VSS.n3197 1.1255
R4270 VSS.n3347 VSS.n3346 1.1255
R4271 VSS.n3345 VSS.n3201 1.1255
R4272 VSS.n3344 VSS.n3343 1.1255
R4273 VSS.n3204 VSS.n3203 1.1255
R4274 VSS.n3206 VSS.n53 1.1255
R4275 VSS.n3209 VSS.n54 1.1255
R4276 VSS.n3332 VSS.n3331 1.1255
R4277 VSS.n3330 VSS.n3210 1.1255
R4278 VSS.n3329 VSS.n3328 1.1255
R4279 VSS.n3212 VSS.n3211 1.1255
R4280 VSS.n3322 VSS.n51 1.1255
R4281 VSS.n3321 VSS.n52 1.1255
R4282 VSS.n3320 VSS.n3216 1.1255
R4283 VSS.n3221 VSS.n3215 1.1255
R4284 VSS.n3314 VSS.n3313 1.1255
R4285 VSS.n3312 VSS.n3220 1.1255
R4286 VSS.n3311 VSS.n3310 1.1255
R4287 VSS.n3222 VSS.n49 1.1255
R4288 VSS.n3224 VSS.n50 1.1255
R4289 VSS.n3229 VSS.n3227 1.1255
R4290 VSS.n3299 VSS.n3298 1.1255
R4291 VSS.n3297 VSS.n3228 1.1255
R4292 VSS.n3296 VSS.n3295 1.1255
R4293 VSS.n3230 VSS.n47 1.1255
R4294 VSS.n3289 VSS.n48 1.1255
R4295 VSS.n3288 VSS.n3287 1.1255
R4296 VSS.n3286 VSS.n3234 1.1255
R4297 VSS.n3285 VSS.n3284 1.1255
R4298 VSS.n46 VSS.n45 1.1255
R4299 VSS.n3435 VSS.n3434 1.1255
R4300 VSS.n67 VSS.n66 1.1255
R4301 VSS.n3409 VSS.n3406 1.1255
R4302 VSS.n3413 VSS.n3412 1.1255
R4303 VSS.n3414 VSS.n3405 1.1255
R4304 VSS.n3416 VSS.n3415 1.1255
R4305 VSS.n3404 VSS.n3403 1.1255
R4306 VSS.n3421 VSS.n3420 1.1255
R4307 VSS.n3170 VSS.n3168 1.1255
R4308 VSS.n3426 VSS.n3425 1.1255
R4309 VSS.n3401 VSS.n3169 1.1255
R4310 VSS.n3400 VSS.n3399 1.1255
R4311 VSS.n3397 VSS.n3171 1.1255
R4312 VSS.n3175 VSS.n3172 1.1255
R4313 VSS.n3393 VSS.n3392 1.1255
R4314 VSS.n3176 VSS.n3174 1.1255
R4315 VSS.n3388 VSS.n3387 1.1255
R4316 VSS.n3180 VSS.n3179 1.1255
R4317 VSS.n3383 VSS.n3382 1.1255
R4318 VSS.n3381 VSS.n3182 1.1255
R4319 VSS.n3186 VSS.n3183 1.1255
R4320 VSS.n3377 VSS.n3376 1.1255
R4321 VSS.n3372 VSS.n3185 1.1255
R4322 VSS.n3371 VSS.n3188 1.1255
R4323 VSS.n3191 VSS.n3187 1.1255
R4324 VSS.n3367 VSS.n3366 1.1255
R4325 VSS.n3192 VSS.n3190 1.1255
R4326 VSS.n3362 VSS.n3361 1.1255
R4327 VSS.n3195 VSS.n3194 1.1255
R4328 VSS.n3357 VSS.n3356 1.1255
R4329 VSS.n3354 VSS.n3196 1.1255
R4330 VSS.n3353 VSS.n3352 1.1255
R4331 VSS.n3198 VSS.n3197 1.1255
R4332 VSS.n3348 VSS.n3347 1.1255
R4333 VSS.n3201 VSS.n3200 1.1255
R4334 VSS.n3343 VSS.n3342 1.1255
R4335 VSS.n3338 VSS.n3204 1.1255
R4336 VSS.n3337 VSS.n3206 1.1255
R4337 VSS.n3209 VSS.n3205 1.1255
R4338 VSS.n3333 VSS.n3332 1.1255
R4339 VSS.n3210 VSS.n3208 1.1255
R4340 VSS.n3328 VSS.n3327 1.1255
R4341 VSS.n3213 VSS.n3212 1.1255
R4342 VSS.n3323 VSS.n3322 1.1255
R4343 VSS.n3321 VSS.n3214 1.1255
R4344 VSS.n3320 VSS.n3319 1.1255
R4345 VSS.n3217 VSS.n3215 1.1255
R4346 VSS.n3315 VSS.n3314 1.1255
R4347 VSS.n3220 VSS.n3219 1.1255
R4348 VSS.n3310 VSS.n3309 1.1255
R4349 VSS.n3305 VSS.n3222 1.1255
R4350 VSS.n3304 VSS.n3224 1.1255
R4351 VSS.n3227 VSS.n3223 1.1255
R4352 VSS.n3300 VSS.n3299 1.1255
R4353 VSS.n3228 VSS.n3226 1.1255
R4354 VSS.n3295 VSS.n3294 1.1255
R4355 VSS.n3231 VSS.n3230 1.1255
R4356 VSS.n3290 VSS.n3289 1.1255
R4357 VSS.n3288 VSS.n3233 1.1255
R4358 VSS.n3235 VSS.n3234 1.1255
R4359 VSS.n3284 VSS.n3283 1.1255
R4360 VSS.n3279 VSS.n45 1.1255
R4361 VSS.n3434 VSS.n3433 1.1255
R4362 VSS.n3281 VSS.n3279 1.1255
R4363 VSS.n3283 VSS.n3282 1.1255
R4364 VSS.n3280 VSS.n3235 1.1255
R4365 VSS.n3233 VSS.n3232 1.1255
R4366 VSS.n3291 VSS.n3290 1.1255
R4367 VSS.n3292 VSS.n3231 1.1255
R4368 VSS.n3294 VSS.n3293 1.1255
R4369 VSS.n3226 VSS.n3225 1.1255
R4370 VSS.n3301 VSS.n3300 1.1255
R4371 VSS.n3302 VSS.n3223 1.1255
R4372 VSS.n3304 VSS.n3303 1.1255
R4373 VSS.n3307 VSS.n3305 1.1255
R4374 VSS.n3309 VSS.n3308 1.1255
R4375 VSS.n3306 VSS.n3219 1.1255
R4376 VSS.n3316 VSS.n3315 1.1255
R4377 VSS.n3317 VSS.n3217 1.1255
R4378 VSS.n3319 VSS.n3318 1.1255
R4379 VSS.n3218 VSS.n3214 1.1255
R4380 VSS.n3324 VSS.n3323 1.1255
R4381 VSS.n3325 VSS.n3213 1.1255
R4382 VSS.n3327 VSS.n3326 1.1255
R4383 VSS.n3208 VSS.n3207 1.1255
R4384 VSS.n3334 VSS.n3333 1.1255
R4385 VSS.n3335 VSS.n3205 1.1255
R4386 VSS.n3337 VSS.n3336 1.1255
R4387 VSS.n3340 VSS.n3338 1.1255
R4388 VSS.n3342 VSS.n3341 1.1255
R4389 VSS.n3339 VSS.n3200 1.1255
R4390 VSS.n3349 VSS.n3348 1.1255
R4391 VSS.n3350 VSS.n3198 1.1255
R4392 VSS.n3352 VSS.n3351 1.1255
R4393 VSS.n3199 VSS.n3196 1.1255
R4394 VSS.n3358 VSS.n3357 1.1255
R4395 VSS.n3359 VSS.n3195 1.1255
R4396 VSS.n3361 VSS.n3360 1.1255
R4397 VSS.n3190 VSS.n3189 1.1255
R4398 VSS.n3368 VSS.n3367 1.1255
R4399 VSS.n3369 VSS.n3187 1.1255
R4400 VSS.n3371 VSS.n3370 1.1255
R4401 VSS.n3374 VSS.n3372 1.1255
R4402 VSS.n3376 VSS.n3375 1.1255
R4403 VSS.n3373 VSS.n3186 1.1255
R4404 VSS.n3182 VSS.n3181 1.1255
R4405 VSS.n3384 VSS.n3383 1.1255
R4406 VSS.n3385 VSS.n3180 1.1255
R4407 VSS.n3387 VSS.n3386 1.1255
R4408 VSS.n3174 VSS.n3173 1.1255
R4409 VSS.n3394 VSS.n3393 1.1255
R4410 VSS.n3395 VSS.n3172 1.1255
R4411 VSS.n3397 VSS.n3396 1.1255
R4412 VSS.n3399 VSS.n3398 1.1255
R4413 VSS.n3169 VSS.n3167 1.1255
R4414 VSS.n3427 VSS.n3426 1.1255
R4415 VSS.n3168 VSS.n3166 1.1255
R4416 VSS.n3420 VSS.n3419 1.1255
R4417 VSS.n3418 VSS.n3404 1.1255
R4418 VSS.n3417 VSS.n3416 1.1255
R4419 VSS.n3410 VSS.n3405 1.1255
R4420 VSS.n3412 VSS.n3411 1.1255
R4421 VSS.n3409 VSS.n69 1.1255
R4422 VSS.n3431 VSS.n67 1.1255
R4423 VSS.n3433 VSS.n3432 1.1255
R4424 VSS.n1413 VSS.n1082 1.0535
R4425 VSS.n1759 VSS.n1758 1.05237
R4426 VSS.n1356 VSS.n1079 0.977
R4427 VSS.n14 VSS.n0 0.94832
R4428 VSS.n1886 VSS.n433 0.939203
R4429 VSS.n1889 VSS.n433 0.939203
R4430 VSS.n1946 VSS.n311 0.939203
R4431 VSS.n1913 VSS.n311 0.939203
R4432 VSS.n326 VSS.n325 0.939203
R4433 VSS.n325 VSS.n324 0.939203
R4434 VSS.n1806 VSS.n553 0.939203
R4435 VSS.n1808 VSS.n553 0.939203
R4436 VSS.n1790 VSS.n555 0.939203
R4437 VSS.n1778 VSS.n555 0.939203
R4438 VSS.n1797 VSS.n555 0.939203
R4439 VSS.n1800 VSS.n555 0.939203
R4440 VSS.n1870 VSS.n435 0.939203
R4441 VSS.n1858 VSS.n435 0.939203
R4442 VSS.n1877 VSS.n435 0.939203
R4443 VSS.n1880 VSS.n435 0.939203
R4444 VSS.n1930 VSS.n313 0.939203
R4445 VSS.n1919 VSS.n313 0.939203
R4446 VSS.n1937 VSS.n313 0.939203
R4447 VSS.n1940 VSS.n313 0.939203
R4448 VSS.n353 VSS.n314 0.939203
R4449 VSS.n353 VSS.n315 0.939203
R4450 VSS.n353 VSS.n316 0.939203
R4451 VSS.n353 VSS.n317 0.939203
R4452 VSS.n3042 VSS.n3041 0.939203
R4453 VSS.n3041 VSS.n170 0.939203
R4454 VSS.n3041 VSS.n169 0.939203
R4455 VSS.n3041 VSS.n168 0.939203
R4456 VSS.n2879 VSS.n2878 0.939203
R4457 VSS.n2879 VSS.n268 0.939203
R4458 VSS.n384 VSS.n378 0.939203
R4459 VSS.n387 VSS.n378 0.939203
R4460 VSS.n2606 VSS.n2605 0.939203
R4461 VSS.n2606 VSS.n415 0.939203
R4462 VSS.n504 VSS.n496 0.939203
R4463 VSS.n507 VSS.n496 0.939203
R4464 VSS.n2339 VSS.n2338 0.939203
R4465 VSS.n2339 VSS.n535 0.939203
R4466 VSS.n2841 VSS.n2840 0.939203
R4467 VSS.n2841 VSS.n288 0.939203
R4468 VSS.n2745 VSS.n2744 0.939203
R4469 VSS.n2745 VSS.n358 0.939203
R4470 VSS.n444 VSS.n432 0.939203
R4471 VSS.n440 VSS.n432 0.939203
R4472 VSS.n2470 VSS.n478 0.939203
R4473 VSS.n2470 VSS.n2469 0.939203
R4474 VSS.n565 VSS.n552 0.939203
R4475 VSS.n561 VSS.n552 0.939203
R4476 VSS.n1783 VSS.n552 0.939203
R4477 VSS.n1781 VSS.n552 0.939203
R4478 VSS.n1863 VSS.n432 0.939203
R4479 VSS.n1861 VSS.n432 0.939203
R4480 VSS.n2745 VSS.n357 0.939203
R4481 VSS.n2745 VSS.n356 0.939203
R4482 VSS.n2841 VSS.n287 0.939203
R4483 VSS.n2841 VSS.n286 0.939203
R4484 VSS.n2470 VSS.n475 0.939203
R4485 VSS.n2470 VSS.n473 0.939203
R4486 VSS.n2074 VSS.n556 0.939203
R4487 VSS.n2065 VSS.n556 0.939203
R4488 VSS.n2081 VSS.n556 0.939203
R4489 VSS.n2084 VSS.n556 0.939203
R4490 VSS.n2091 VSS.n2090 0.939203
R4491 VSS.n2091 VSS.n2053 0.939203
R4492 VSS.n714 VSS.n129 0.939203
R4493 VSS.n712 VSS.n129 0.939203
R4494 VSS.n721 VSS.n117 0.939203
R4495 VSS.n709 VSS.n117 0.939203
R4496 VSS.n728 VSS.n117 0.939203
R4497 VSS.n731 VSS.n117 0.939203
R4498 VSS.n737 VSS.n700 0.939203
R4499 VSS.n740 VSS.n700 0.939203
R4500 VSS.n215 VSS.n129 0.939203
R4501 VSS.n220 VSS.n129 0.939203
R4502 VSS.n2920 VSS.n244 0.939203
R4503 VSS.n2923 VSS.n244 0.939203
R4504 VSS.n810 VSS.n151 0.939203
R4505 VSS.n804 VSS.n151 0.939203
R4506 VSS.n802 VSS.n151 0.939203
R4507 VSS.n895 VSS.n789 0.939203
R4508 VSS.n829 VSS.n151 0.939203
R4509 VSS.n815 VSS.n151 0.939203
R4510 VSS.n822 VSS.n151 0.939203
R4511 VSS.n817 VSS.n151 0.939203
R4512 VSS.n846 VSS.n19 0.939203
R4513 VSS.n856 VSS.n19 0.939203
R4514 VSS.n844 VSS.n19 0.939203
R4515 VSS.n3082 VSS.n133 0.939203
R4516 VSS.n3085 VSS.n133 0.939203
R4517 VSS.n757 VSS.n81 0.939203
R4518 VSS.n760 VSS.n81 0.939203
R4519 VSS.n767 VSS.n80 0.939203
R4520 VSS.n773 VSS.n80 0.939203
R4521 VSS.n775 VSS.n80 0.939203
R4522 VSS.n781 VSS.n80 0.939203
R4523 VSS.n908 VSS.n80 0.939203
R4524 VSS.n914 VSS.n80 0.939203
R4525 VSS.n916 VSS.n80 0.939203
R4526 VSS.n922 VSS.n80 0.939203
R4527 VSS.n924 VSS.n80 0.939203
R4528 VSS.n930 VSS.n80 0.939203
R4529 VSS.n932 VSS.n80 0.939203
R4530 VSS.n938 VSS.n80 0.939203
R4531 VSS.n940 VSS.n80 0.939203
R4532 VSS.n1496 VSS.n1407 0.93088
R4533 VSS.n1631 VSS.n1629 0.9185
R4534 VSS.n195 VSS.n194 0.915775
R4535 VSS.n3449 VSS.n3448 0.907605
R4536 VSS.n615 VSS.n612 0.904493
R4537 VSS.n3278 VSS.n3277 0.9005
R4538 VSS.n3463 VSS.n14 0.871619
R4539 VSS.n1403 VSS.n1105 0.867167
R4540 VSS.n1404 VSS.n1403 0.867167
R4541 VSS.n31 VSS.n30 0.867167
R4542 VSS.n3455 VSS.n3454 0.867167
R4543 VSS.n3454 VSS.n3453 0.867167
R4544 VSS.n963 VSS.t338 0.833115
R4545 VSS.n163 VSS.t89 0.8195
R4546 VSS.n163 VSS.t193 0.8195
R4547 VSS.n164 VSS.t5 0.8195
R4548 VSS.n164 VSS.t143 0.8195
R4549 VSS.n1592 VSS.n1591 0.807125
R4550 VSS.n1365 VSS.n1364 0.779896
R4551 VSS.n850 VSS.n848 0.77784
R4552 VSS.t189 VSS.n3435 0.758022
R4553 VSS.n29 VSS.n28 0.73471
R4554 VSS.n1200 VSS.n1161 0.705167
R4555 VSS.n1166 VSS.n1161 0.705167
R4556 VSS.n1193 VSS.n1161 0.705167
R4557 VSS.n1187 VSS.n1161 0.705167
R4558 VSS.n1185 VSS.n1161 0.705167
R4559 VSS.n1179 VSS.n1161 0.705167
R4560 VSS.n1177 VSS.n1161 0.705167
R4561 VSS.n1172 VSS.n1161 0.705167
R4562 VSS.n1344 VSS.n1229 0.705167
R4563 VSS.n1344 VSS.n1230 0.705167
R4564 VSS.n1344 VSS.n1231 0.705167
R4565 VSS.n1344 VSS.n1232 0.705167
R4566 VSS.n1344 VSS.n1233 0.705167
R4567 VSS.n1344 VSS.n1234 0.705167
R4568 VSS.n1344 VSS.n1235 0.705167
R4569 VSS.n1344 VSS.n1236 0.705167
R4570 VSS.n1690 VSS.n1064 0.698475
R4571 VSS.n1690 VSS.n1065 0.698475
R4572 VSS.n1690 VSS.n1066 0.698475
R4573 VSS.n1690 VSS.n1067 0.698475
R4574 VSS.n1690 VSS.n1068 0.698475
R4575 VSS.n1690 VSS.n1069 0.698475
R4576 VSS.n1690 VSS.n1689 0.698475
R4577 VSS.n1536 VSS.n1513 0.660831
R4578 VSS.n2361 VSS.n2360 0.660831
R4579 VSS.n2417 VSS.n2394 0.660831
R4580 VSS.n2628 VSS.n2627 0.660831
R4581 VSS.n2689 VSS.n2661 0.660831
R4582 VSS.n2900 VSS.n255 0.660831
R4583 VSS.n3440 VSS.n45 0.64962
R4584 VSS.n2131 VSS.n2130 0.642811
R4585 VSS.n1147 VSS.n1109 0.608375
R4586 VSS.n1568 VSS.n1567 0.608
R4587 VSS.n1758 VSS.n620 0.58325
R4588 VSS.n944 VSS.n41 0.567737
R4589 VSS.n852 VSS.n22 0.553526
R4590 VSS.n1661 VSS.n1071 0.545237
R4591 VSS.n1690 VSS.n1063 0.538771
R4592 VSS.n1590 VSS.n1416 0.532146
R4593 VSS.n1662 VSS.n1661 0.513263
R4594 VSS.n1695 VSS.n1694 0.50099
R4595 VSS.n1754 VSS.n1753 0.5005
R4596 VSS.n1721 VSS.n1024 0.5005
R4597 VSS.n1717 VSS.n1019 0.5005
R4598 VSS.n1723 VSS.n1027 0.5005
R4599 VSS.n1714 VSS.n1018 0.5005
R4600 VSS.n1725 VSS.n1030 0.5005
R4601 VSS.n1713 VSS.n1017 0.5005
R4602 VSS.n1727 VSS.n1033 0.5005
R4603 VSS.n1712 VSS.n1016 0.5005
R4604 VSS.n1729 VSS.n1036 0.5005
R4605 VSS.n1711 VSS.n1015 0.5005
R4606 VSS.n1731 VSS.n1039 0.5005
R4607 VSS.n1710 VSS.n1014 0.5005
R4608 VSS.n1733 VSS.n1042 0.5005
R4609 VSS.n1709 VSS.n1013 0.5005
R4610 VSS.n1735 VSS.n1044 0.5005
R4611 VSS.n1708 VSS.n1707 0.5005
R4612 VSS.n1748 VSS.n1045 0.5005
R4613 VSS.n1702 VSS.n1050 0.5005
R4614 VSS.n1751 VSS.n1750 0.5005
R4615 VSS.n1021 VSS.n622 0.5005
R4616 VSS.n1756 VSS.n627 0.5005
R4617 VSS.n1312 VSS.n1261 0.476553
R4618 VSS.n1342 VSS.n1225 0.471816
R4619 VSS.n1696 VSS.n1054 0.460063
R4620 VSS.n1394 VSS.n1105 0.458789
R4621 VSS.n1609 VSS.n1105 0.458789
R4622 VSS.n3456 VSS.n3455 0.458789
R4623 VSS.n3455 VSS.n23 0.458789
R4624 VSS.n3275 VSS.n3236 0.452273
R4625 VSS.n1213 VSS.n1212 0.43349
R4626 VSS.n1204 VSS.n1203 0.419711
R4627 VSS.n30 VSS.n12 0.413789
R4628 VSS.n1380 VSS.n1379 0.4082
R4629 VSS.n1356 VSS.n614 0.4005
R4630 VSS.n614 VSS.n603 0.4005
R4631 VSS.n8 VSS.n1 0.394162
R4632 VSS.n1215 VSS.n1056 0.39128
R4633 VSS.n1203 VSS.n1155 0.3866
R4634 VSS.n1386 VSS.n1385 0.3668
R4635 VSS.n1687 VSS.n1058 0.365237
R4636 VSS.n1687 VSS.n1686 0.365237
R4637 VSS.n1686 VSS.n1685 0.365237
R4638 VSS.n1685 VSS.n1682 0.365237
R4639 VSS.n1682 VSS.n1681 0.365237
R4640 VSS.n1681 VSS.n1678 0.365237
R4641 VSS.n1678 VSS.n1677 0.365237
R4642 VSS.n1677 VSS.n1674 0.365237
R4643 VSS.n1674 VSS.n1673 0.365237
R4644 VSS.n1673 VSS.n1670 0.365237
R4645 VSS.n1670 VSS.n1669 0.365237
R4646 VSS.n1669 VSS.n1666 0.365237
R4647 VSS.n1666 VSS.n1665 0.365237
R4648 VSS.n1665 VSS.n1662 0.365237
R4649 VSS.n1342 VSS.n1341 0.3605
R4650 VSS.n1341 VSS.n1340 0.3605
R4651 VSS.n1340 VSS.n1337 0.3605
R4652 VSS.n1337 VSS.n1336 0.3605
R4653 VSS.n1336 VSS.n1333 0.3605
R4654 VSS.n1333 VSS.n1332 0.3605
R4655 VSS.n1332 VSS.n1329 0.3605
R4656 VSS.n1329 VSS.n1328 0.3605
R4657 VSS.n1328 VSS.n1325 0.3605
R4658 VSS.n1325 VSS.n1324 0.3605
R4659 VSS.n1324 VSS.n1321 0.3605
R4660 VSS.n1321 VSS.n1320 0.3605
R4661 VSS.n1320 VSS.n1317 0.3605
R4662 VSS.n1317 VSS.n1316 0.3605
R4663 VSS.n1316 VSS.n1313 0.3605
R4664 VSS.n1313 VSS.n1312 0.3605
R4665 VSS.n1383 VSS.n1154 0.3605
R4666 VSS.n1383 VSS.n1382 0.3605
R4667 VSS.n1382 VSS.n1155 0.3605
R4668 VSS.n1202 VSS.n1165 0.3605
R4669 VSS.n1197 VSS.n1165 0.3605
R4670 VSS.n1197 VSS.n1196 0.3605
R4671 VSS.n1196 VSS.n1167 0.3605
R4672 VSS.n1191 VSS.n1167 0.3605
R4673 VSS.n1191 VSS.n1190 0.3605
R4674 VSS.n1190 VSS.n1189 0.3605
R4675 VSS.n1189 VSS.n1169 0.3605
R4676 VSS.n1183 VSS.n1169 0.3605
R4677 VSS.n1183 VSS.n1182 0.3605
R4678 VSS.n1182 VSS.n1181 0.3605
R4679 VSS.n1181 VSS.n1171 0.3605
R4680 VSS.n1175 VSS.n1171 0.3605
R4681 VSS.n1175 VSS.n1174 0.3605
R4682 VSS.n1174 VSS.n1156 0.3605
R4683 VSS.n1385 VSS.n1152 0.3578
R4684 VSS.n1394 VSS.n1393 0.355763
R4685 VSS.n1380 VSS.n1152 0.3461
R4686 VSS.n1635 VSS.n1634 0.3317
R4687 VSS.n1634 VSS.n1080 0.3317
R4688 VSS.n1648 VSS.n1647 0.3317
R4689 VSS.n1393 VSS.n1392 0.3255
R4690 VSS.n1148 VSS.n1095 0.32075
R4691 VSS.n1373 VSS.n1372 0.313132
R4692 VSS.n1372 VSS.n1371 0.313132
R4693 VSS.n1371 VSS.n1205 0.313132
R4694 VSS.n1349 VSS.n1224 0.313132
R4695 VSS.n1349 VSS.n1348 0.313132
R4696 VSS.n1348 VSS.n1347 0.313132
R4697 VSS.n1288 VSS.n1264 0.313132
R4698 VSS.n1288 VSS.n1287 0.313132
R4699 VSS.n1287 VSS.n1286 0.313132
R4700 VSS.n1286 VSS.n1265 0.313132
R4701 VSS.n1280 VSS.n1265 0.313132
R4702 VSS.n1280 VSS.n1279 0.313132
R4703 VSS.n1279 VSS.n1278 0.313132
R4704 VSS.n1278 VSS.n1270 0.313132
R4705 VSS.n1272 VSS.n1270 0.313132
R4706 VSS.n1272 VSS.n1271 0.313132
R4707 VSS.n1377 VSS.n1158 0.313132
R4708 VSS.n1238 VSS.n1158 0.313132
R4709 VSS.n1239 VSS.n1238 0.313132
R4710 VSS.n1240 VSS.n1239 0.313132
R4711 VSS.n1254 VSS.n1240 0.313132
R4712 VSS.n1255 VSS.n1254 0.313132
R4713 VSS.n1256 VSS.n1255 0.313132
R4714 VSS.n1257 VSS.n1256 0.313132
R4715 VSS.n1259 VSS.n1257 0.313132
R4716 VSS.n1260 VSS.n1259 0.313132
R4717 VSS.n1308 VSS.n1307 0.313132
R4718 VSS.n1307 VSS.n1306 0.313132
R4719 VSS.n1306 VSS.n1292 0.313132
R4720 VSS.n1300 VSS.n1292 0.313132
R4721 VSS.n1300 VSS.n1299 0.313132
R4722 VSS.n1299 VSS.n1298 0.313132
R4723 VSS.n1298 VSS.n1073 0.313132
R4724 VSS.n1656 VSS.n1073 0.313132
R4725 VSS.n1657 VSS.n1656 0.313132
R4726 VSS.n1658 VSS.n1657 0.313132
R4727 VSS.n1692 VSS.n1058 0.311947
R4728 VSS.n1216 VSS.n1205 0.311947
R4729 VSS.n1378 VSS.n1157 0.310763
R4730 VSS.n1357 VSS.n1071 0.310763
R4731 VSS.n1620 VSS.n1096 0.305
R4732 VSS.n1358 VSS.n1357 0.3015
R4733 VSS.n1203 VSS.n1202 0.294184
R4734 VSS.n1109 VSS.n1091 0.289389
R4735 VSS.n1624 VSS.n1091 0.289389
R4736 VSS.n1642 VSS.n1641 0.289389
R4737 VSS.n1641 VSS.n1062 0.289389
R4738 VSS.n1148 VSS.n1147 0.28775
R4739 VSS.n1582 VSS.n1581 0.286527
R4740 VSS.n1581 VSS.n1580 0.286527
R4741 VSS.n1213 VSS.n1154 0.2849
R4742 VSS.n1214 VSS.n1213 0.27473
R4743 VSS.n847 VSS.n20 0.27425
R4744 VSS.n1212 VSS.n1151 0.2741
R4745 VSS.n1224 VSS.n1216 0.2705
R4746 VSS.n1387 VSS.n1150 0.2705
R4747 VSS.n1591 VSS.n1414 0.269375
R4748 VSS.n3157 VSS.n82 0.265655
R4749 VSS.n1054 VSS.n619 0.254021
R4750 VSS.n616 VSS.n601 0.254021
R4751 VSS.n2177 VSS.n601 0.254021
R4752 VSS.n2178 VSS.n2177 0.254021
R4753 VSS.n2178 VSS.n599 0.254021
R4754 VSS.n2182 VSS.n599 0.254021
R4755 VSS.n2183 VSS.n2182 0.254021
R4756 VSS.n2183 VSS.n596 0.254021
R4757 VSS.n2203 VSS.n2187 0.254021
R4758 VSS.n2203 VSS.n2202 0.254021
R4759 VSS.n2202 VSS.n2201 0.254021
R4760 VSS.n2201 VSS.n2189 0.254021
R4761 VSS.n2196 VSS.n2189 0.254021
R4762 VSS.n2196 VSS.n2195 0.254021
R4763 VSS.n2195 VSS.n2194 0.254021
R4764 VSS.n1466 VSS.n1465 0.254021
R4765 VSS.n1467 VSS.n1466 0.254021
R4766 VSS.n1468 VSS.n1467 0.254021
R4767 VSS.n1472 VSS.n1468 0.254021
R4768 VSS.n1473 VSS.n1472 0.254021
R4769 VSS.n1474 VSS.n1473 0.254021
R4770 VSS.n1474 VSS.n1459 0.254021
R4771 VSS.n1481 VSS.n1459 0.254021
R4772 VSS.n1482 VSS.n1481 0.254021
R4773 VSS.n1483 VSS.n1482 0.254021
R4774 VSS.n1487 VSS.n1486 0.254021
R4775 VSS.n1488 VSS.n1487 0.254021
R4776 VSS.n1488 VSS.n1454 0.254021
R4777 VSS.n1494 VSS.n1454 0.254021
R4778 VSS.n1495 VSS.n1494 0.254021
R4779 VSS.n1503 VSS.n1495 0.254021
R4780 VSS.n1503 VSS.n1502 0.254021
R4781 VSS.n1502 VSS.n1501 0.254021
R4782 VSS.n1501 VSS.n1498 0.254021
R4783 VSS.n1498 VSS.n1497 0.254021
R4784 VSS.n1355 VSS.n1354 0.248119
R4785 VSS.n1355 VSS.n1090 0.248119
R4786 VSS.n36 VSS.n35 0.248119
R4787 VSS.t332 VSS.n36 0.248119
R4788 VSS.n1421 VSS.n1095 0.243993
R4789 VSS.n1569 VSS.n1568 0.243993
R4790 VSS.n1626 VSS.n1089 0.2408
R4791 VSS.n2151 VSS.n615 0.238393
R4792 VSS.n217 VSS.n123 0.237342
R4793 VSS.n218 VSS.n217 0.237342
R4794 VSS.n218 VSS.n213 0.237342
R4795 VSS.n213 VSS.n212 0.237342
R4796 VSS.n226 VSS.n212 0.237342
R4797 VSS.n227 VSS.n226 0.237342
R4798 VSS.n228 VSS.n227 0.237342
R4799 VSS.n228 VSS.n208 0.237342
R4800 VSS.n234 VSS.n208 0.237342
R4801 VSS.n235 VSS.n234 0.237342
R4802 VSS.n2957 VSS.n235 0.237342
R4803 VSS.n2957 VSS.n2956 0.237342
R4804 VSS.n2956 VSS.n2955 0.237342
R4805 VSS.n2955 VSS.n236 0.237342
R4806 VSS.n2949 VSS.n236 0.237342
R4807 VSS.n2949 VSS.n2948 0.237342
R4808 VSS.n2948 VSS.n2947 0.237342
R4809 VSS.n2947 VSS.n240 0.237342
R4810 VSS.n2919 VSS.n240 0.237342
R4811 VSS.n2919 VSS.n2918 0.237342
R4812 VSS.n2925 VSS.n2918 0.237342
R4813 VSS.n742 VSS.n702 0.237342
R4814 VSS.n703 VSS.n702 0.237342
R4815 VSS.n735 VSS.n703 0.237342
R4816 VSS.n735 VSS.n734 0.237342
R4817 VSS.n734 VSS.n733 0.237342
R4818 VSS.n733 VSS.n705 0.237342
R4819 VSS.n706 VSS.n705 0.237342
R4820 VSS.n726 VSS.n706 0.237342
R4821 VSS.n726 VSS.n725 0.237342
R4822 VSS.n725 VSS.n724 0.237342
R4823 VSS.n724 VSS.n708 0.237342
R4824 VSS.n719 VSS.n708 0.237342
R4825 VSS.n719 VSS.n718 0.237342
R4826 VSS.n718 VSS.n717 0.237342
R4827 VSS.n717 VSS.n711 0.237342
R4828 VSS.n711 VSS.n124 0.237342
R4829 VSS.n175 VSS.n162 0.237342
R4830 VSS.n176 VSS.n175 0.237342
R4831 VSS.n179 VSS.n176 0.237342
R4832 VSS.n180 VSS.n179 0.237342
R4833 VSS.n183 VSS.n180 0.237342
R4834 VSS.n185 VSS.n183 0.237342
R4835 VSS.n567 VSS.n560 0.237342
R4836 VSS.n562 VSS.n560 0.237342
R4837 VSS.n562 VSS.n550 0.237342
R4838 VSS.n2306 VSS.n550 0.237342
R4839 VSS.n2307 VSS.n2306 0.237342
R4840 VSS.n2308 VSS.n2307 0.237342
R4841 VSS.n2308 VSS.n546 0.237342
R4842 VSS.n2314 VSS.n546 0.237342
R4843 VSS.n2315 VSS.n2314 0.237342
R4844 VSS.n2316 VSS.n2315 0.237342
R4845 VSS.n2316 VSS.n542 0.237342
R4846 VSS.n2322 VSS.n542 0.237342
R4847 VSS.n2323 VSS.n2322 0.237342
R4848 VSS.n2324 VSS.n2323 0.237342
R4849 VSS.n2324 VSS.n538 0.237342
R4850 VSS.n2331 VSS.n538 0.237342
R4851 VSS.n2332 VSS.n2331 0.237342
R4852 VSS.n2336 VSS.n2332 0.237342
R4853 VSS.n2336 VSS.n2335 0.237342
R4854 VSS.n2335 VSS.n2334 0.237342
R4855 VSS.n2334 VSS.n530 0.237342
R4856 VSS.n481 VSS.n468 0.237342
R4857 VSS.n2467 VSS.n481 0.237342
R4858 VSS.n2467 VSS.n2466 0.237342
R4859 VSS.n2466 VSS.n2465 0.237342
R4860 VSS.n2465 VSS.n482 0.237342
R4861 VSS.n2459 VSS.n482 0.237342
R4862 VSS.n2459 VSS.n2458 0.237342
R4863 VSS.n2458 VSS.n2457 0.237342
R4864 VSS.n2457 VSS.n486 0.237342
R4865 VSS.n2451 VSS.n486 0.237342
R4866 VSS.n2451 VSS.n2450 0.237342
R4867 VSS.n2450 VSS.n2449 0.237342
R4868 VSS.n2449 VSS.n490 0.237342
R4869 VSS.n2443 VSS.n490 0.237342
R4870 VSS.n2443 VSS.n2442 0.237342
R4871 VSS.n2442 VSS.n2441 0.237342
R4872 VSS.n2441 VSS.n494 0.237342
R4873 VSS.n502 VSS.n494 0.237342
R4874 VSS.n502 VSS.n501 0.237342
R4875 VSS.n501 VSS.n500 0.237342
R4876 VSS.n509 VSS.n500 0.237342
R4877 VSS.n446 VSS.n439 0.237342
R4878 VSS.n441 VSS.n439 0.237342
R4879 VSS.n441 VSS.n430 0.237342
R4880 VSS.n2573 VSS.n430 0.237342
R4881 VSS.n2574 VSS.n2573 0.237342
R4882 VSS.n2575 VSS.n2574 0.237342
R4883 VSS.n2575 VSS.n426 0.237342
R4884 VSS.n2581 VSS.n426 0.237342
R4885 VSS.n2582 VSS.n2581 0.237342
R4886 VSS.n2583 VSS.n2582 0.237342
R4887 VSS.n2583 VSS.n422 0.237342
R4888 VSS.n2589 VSS.n422 0.237342
R4889 VSS.n2590 VSS.n2589 0.237342
R4890 VSS.n2591 VSS.n2590 0.237342
R4891 VSS.n2591 VSS.n418 0.237342
R4892 VSS.n2598 VSS.n418 0.237342
R4893 VSS.n2599 VSS.n2598 0.237342
R4894 VSS.n2603 VSS.n2599 0.237342
R4895 VSS.n2603 VSS.n2602 0.237342
R4896 VSS.n2602 VSS.n2601 0.237342
R4897 VSS.n2601 VSS.n410 0.237342
R4898 VSS.n2742 VSS.n2741 0.237342
R4899 VSS.n2741 VSS.n2740 0.237342
R4900 VSS.n2740 VSS.n2738 0.237342
R4901 VSS.n2738 VSS.n362 0.237342
R4902 VSS.n364 VSS.n362 0.237342
R4903 VSS.n367 VSS.n364 0.237342
R4904 VSS.n2730 VSS.n367 0.237342
R4905 VSS.n2730 VSS.n2729 0.237342
R4906 VSS.n2729 VSS.n2728 0.237342
R4907 VSS.n2728 VSS.n368 0.237342
R4908 VSS.n2722 VSS.n368 0.237342
R4909 VSS.n2722 VSS.n2721 0.237342
R4910 VSS.n2721 VSS.n2720 0.237342
R4911 VSS.n2720 VSS.n372 0.237342
R4912 VSS.n2714 VSS.n372 0.237342
R4913 VSS.n2714 VSS.n2713 0.237342
R4914 VSS.n2713 VSS.n2712 0.237342
R4915 VSS.n2712 VSS.n376 0.237342
R4916 VSS.n383 VSS.n376 0.237342
R4917 VSS.n383 VSS.n382 0.237342
R4918 VSS.n389 VSS.n382 0.237342
R4919 VSS.n2838 VSS.n2837 0.237342
R4920 VSS.n2837 VSS.n2836 0.237342
R4921 VSS.n2836 VSS.n283 0.237342
R4922 VSS.n2845 VSS.n283 0.237342
R4923 VSS.n2846 VSS.n2845 0.237342
R4924 VSS.n2847 VSS.n2846 0.237342
R4925 VSS.n2847 VSS.n279 0.237342
R4926 VSS.n2853 VSS.n279 0.237342
R4927 VSS.n2854 VSS.n2853 0.237342
R4928 VSS.n2855 VSS.n2854 0.237342
R4929 VSS.n2855 VSS.n275 0.237342
R4930 VSS.n2861 VSS.n275 0.237342
R4931 VSS.n2862 VSS.n2861 0.237342
R4932 VSS.n2863 VSS.n2862 0.237342
R4933 VSS.n2863 VSS.n271 0.237342
R4934 VSS.n2869 VSS.n271 0.237342
R4935 VSS.n2870 VSS.n2869 0.237342
R4936 VSS.n2876 VSS.n2870 0.237342
R4937 VSS.n2876 VSS.n2875 0.237342
R4938 VSS.n2875 VSS.n2874 0.237342
R4939 VSS.n2874 VSS.n2872 0.237342
R4940 VSS.n320 VSS.n95 0.237342
R4941 VSS.n328 VSS.n320 0.237342
R4942 VSS.n329 VSS.n328 0.237342
R4943 VSS.n351 VSS.n329 0.237342
R4944 VSS.n351 VSS.n350 0.237342
R4945 VSS.n350 VSS.n349 0.237342
R4946 VSS.n349 VSS.n346 0.237342
R4947 VSS.n346 VSS.n345 0.237342
R4948 VSS.n345 VSS.n342 0.237342
R4949 VSS.n342 VSS.n341 0.237342
R4950 VSS.n341 VSS.n338 0.237342
R4951 VSS.n338 VSS.n337 0.237342
R4952 VSS.n337 VSS.n334 0.237342
R4953 VSS.n334 VSS.n333 0.237342
R4954 VSS.n333 VSS.n330 0.237342
R4955 VSS.n330 VSS.n292 0.237342
R4956 VSS.n1950 VSS.n1949 0.237342
R4957 VSS.n1949 VSS.n1912 0.237342
R4958 VSS.n1944 VSS.n1912 0.237342
R4959 VSS.n1944 VSS.n1943 0.237342
R4960 VSS.n1943 VSS.n1942 0.237342
R4961 VSS.n1942 VSS.n1915 0.237342
R4962 VSS.n1916 VSS.n1915 0.237342
R4963 VSS.n1935 VSS.n1916 0.237342
R4964 VSS.n1935 VSS.n1934 0.237342
R4965 VSS.n1934 VSS.n1933 0.237342
R4966 VSS.n1933 VSS.n1918 0.237342
R4967 VSS.n1928 VSS.n1918 0.237342
R4968 VSS.n1928 VSS.n1927 0.237342
R4969 VSS.n1927 VSS.n1926 0.237342
R4970 VSS.n1926 VSS.n1923 0.237342
R4971 VSS.n1923 VSS.n1922 0.237342
R4972 VSS.n1891 VSS.n1851 0.237342
R4973 VSS.n1852 VSS.n1851 0.237342
R4974 VSS.n1884 VSS.n1852 0.237342
R4975 VSS.n1884 VSS.n1883 0.237342
R4976 VSS.n1883 VSS.n1882 0.237342
R4977 VSS.n1882 VSS.n1854 0.237342
R4978 VSS.n1855 VSS.n1854 0.237342
R4979 VSS.n1875 VSS.n1855 0.237342
R4980 VSS.n1875 VSS.n1874 0.237342
R4981 VSS.n1874 VSS.n1873 0.237342
R4982 VSS.n1873 VSS.n1857 0.237342
R4983 VSS.n1868 VSS.n1857 0.237342
R4984 VSS.n1868 VSS.n1867 0.237342
R4985 VSS.n1867 VSS.n1866 0.237342
R4986 VSS.n1866 VSS.n1860 0.237342
R4987 VSS.n1860 VSS.n447 0.237342
R4988 VSS.n1811 VSS.n1810 0.237342
R4989 VSS.n1810 VSS.n1772 0.237342
R4990 VSS.n1804 VSS.n1772 0.237342
R4991 VSS.n1804 VSS.n1803 0.237342
R4992 VSS.n1803 VSS.n1802 0.237342
R4993 VSS.n1802 VSS.n1774 0.237342
R4994 VSS.n1775 VSS.n1774 0.237342
R4995 VSS.n1795 VSS.n1775 0.237342
R4996 VSS.n1795 VSS.n1794 0.237342
R4997 VSS.n1794 VSS.n1793 0.237342
R4998 VSS.n1793 VSS.n1777 0.237342
R4999 VSS.n1788 VSS.n1777 0.237342
R5000 VSS.n1788 VSS.n1787 0.237342
R5001 VSS.n1787 VSS.n1786 0.237342
R5002 VSS.n1786 VSS.n1780 0.237342
R5003 VSS.n1780 VSS.n568 0.237342
R5004 VSS.n2059 VSS.n2057 0.237342
R5005 VSS.n2060 VSS.n2059 0.237342
R5006 VSS.n2088 VSS.n2060 0.237342
R5007 VSS.n2088 VSS.n2087 0.237342
R5008 VSS.n2087 VSS.n2086 0.237342
R5009 VSS.n2086 VSS.n2061 0.237342
R5010 VSS.n2062 VSS.n2061 0.237342
R5011 VSS.n2079 VSS.n2062 0.237342
R5012 VSS.n2079 VSS.n2078 0.237342
R5013 VSS.n2078 VSS.n2077 0.237342
R5014 VSS.n2077 VSS.n2064 0.237342
R5015 VSS.n2072 VSS.n2064 0.237342
R5016 VSS.n2072 VSS.n2071 0.237342
R5017 VSS.n2071 VSS.n2070 0.237342
R5018 VSS.n2070 VSS.n2067 0.237342
R5019 VSS.n2067 VSS.n469 0.237342
R5020 VSS.n787 VSS.n784 0.237342
R5021 VSS.n901 VSS.n787 0.237342
R5022 VSS.n901 VSS.n900 0.237342
R5023 VSS.n900 VSS.n899 0.237342
R5024 VSS.n899 VSS.n788 0.237342
R5025 VSS.n893 VSS.n788 0.237342
R5026 VSS.n893 VSS.n892 0.237342
R5027 VSS.n892 VSS.n891 0.237342
R5028 VSS.n891 VSS.n791 0.237342
R5029 VSS.n800 VSS.n791 0.237342
R5030 VSS.n800 VSS.n799 0.237342
R5031 VSS.n806 VSS.n799 0.237342
R5032 VSS.n807 VSS.n806 0.237342
R5033 VSS.n808 VSS.n807 0.237342
R5034 VSS.n808 VSS.n797 0.237342
R5035 VSS.n813 VSS.n797 0.237342
R5036 VSS.n831 VSS.n814 0.237342
R5037 VSS.n826 VSS.n814 0.237342
R5038 VSS.n826 VSS.n825 0.237342
R5039 VSS.n825 VSS.n816 0.237342
R5040 VSS.n820 VSS.n816 0.237342
R5041 VSS.n820 VSS.n819 0.237342
R5042 VSS.n819 VSS.n155 0.237342
R5043 VSS.n3055 VSS.n155 0.237342
R5044 VSS.n3055 VSS.n3054 0.237342
R5045 VSS.n3054 VSS.n3053 0.237342
R5046 VSS.n3053 VSS.n156 0.237342
R5047 VSS.n3046 VSS.n156 0.237342
R5048 VSS.n3046 VSS.n3045 0.237342
R5049 VSS.n2211 VSS.n585 0.237342
R5050 VSS.n2219 VSS.n585 0.237342
R5051 VSS.n2220 VSS.n2219 0.237342
R5052 VSS.n2221 VSS.n2220 0.237342
R5053 VSS.n2221 VSS.n581 0.237342
R5054 VSS.n2227 VSS.n581 0.237342
R5055 VSS.n2228 VSS.n2227 0.237342
R5056 VSS.n2229 VSS.n2228 0.237342
R5057 VSS.n2229 VSS.n577 0.237342
R5058 VSS.n2235 VSS.n577 0.237342
R5059 VSS.n2236 VSS.n2235 0.237342
R5060 VSS.n2237 VSS.n2236 0.237342
R5061 VSS.n2237 VSS.n573 0.237342
R5062 VSS.n2243 VSS.n573 0.237342
R5063 VSS.n2244 VSS.n2243 0.237342
R5064 VSS.n2245 VSS.n2244 0.237342
R5065 VSS.n2245 VSS.n569 0.237342
R5066 VSS.n2251 VSS.n569 0.237342
R5067 VSS.n2299 VSS.n2298 0.237342
R5068 VSS.n2298 VSS.n2297 0.237342
R5069 VSS.n2297 VSS.n2253 0.237342
R5070 VSS.n2291 VSS.n2253 0.237342
R5071 VSS.n2291 VSS.n2290 0.237342
R5072 VSS.n2290 VSS.n2289 0.237342
R5073 VSS.n2289 VSS.n2257 0.237342
R5074 VSS.n2283 VSS.n2257 0.237342
R5075 VSS.n2283 VSS.n2282 0.237342
R5076 VSS.n2282 VSS.n2281 0.237342
R5077 VSS.n2281 VSS.n2261 0.237342
R5078 VSS.n2275 VSS.n2261 0.237342
R5079 VSS.n2275 VSS.n2274 0.237342
R5080 VSS.n2274 VSS.n2273 0.237342
R5081 VSS.n2273 VSS.n2265 0.237342
R5082 VSS.n2267 VSS.n2265 0.237342
R5083 VSS.n2267 VSS.n470 0.237342
R5084 VSS.n2473 VSS.n470 0.237342
R5085 VSS.n2475 VSS.n464 0.237342
R5086 VSS.n2481 VSS.n464 0.237342
R5087 VSS.n2482 VSS.n2481 0.237342
R5088 VSS.n2483 VSS.n2482 0.237342
R5089 VSS.n2483 VSS.n460 0.237342
R5090 VSS.n2489 VSS.n460 0.237342
R5091 VSS.n2490 VSS.n2489 0.237342
R5092 VSS.n2491 VSS.n2490 0.237342
R5093 VSS.n2491 VSS.n456 0.237342
R5094 VSS.n2497 VSS.n456 0.237342
R5095 VSS.n2498 VSS.n2497 0.237342
R5096 VSS.n2499 VSS.n2498 0.237342
R5097 VSS.n2499 VSS.n452 0.237342
R5098 VSS.n2505 VSS.n452 0.237342
R5099 VSS.n2506 VSS.n2505 0.237342
R5100 VSS.n2507 VSS.n2506 0.237342
R5101 VSS.n2507 VSS.n448 0.237342
R5102 VSS.n2513 VSS.n448 0.237342
R5103 VSS.n2566 VSS.n2565 0.237342
R5104 VSS.n2565 VSS.n2564 0.237342
R5105 VSS.n2564 VSS.n2515 0.237342
R5106 VSS.n2558 VSS.n2515 0.237342
R5107 VSS.n2558 VSS.n2557 0.237342
R5108 VSS.n2557 VSS.n2556 0.237342
R5109 VSS.n2556 VSS.n2519 0.237342
R5110 VSS.n2550 VSS.n2519 0.237342
R5111 VSS.n2550 VSS.n2549 0.237342
R5112 VSS.n2549 VSS.n2548 0.237342
R5113 VSS.n2548 VSS.n2523 0.237342
R5114 VSS.n2542 VSS.n2523 0.237342
R5115 VSS.n2542 VSS.n2541 0.237342
R5116 VSS.n2541 VSS.n2540 0.237342
R5117 VSS.n2540 VSS.n2527 0.237342
R5118 VSS.n2534 VSS.n2527 0.237342
R5119 VSS.n2534 VSS.n2533 0.237342
R5120 VSS.n2533 VSS.n2532 0.237342
R5121 VSS.n2751 VSS.n309 0.237342
R5122 VSS.n2752 VSS.n2751 0.237342
R5123 VSS.n2753 VSS.n2752 0.237342
R5124 VSS.n2753 VSS.n305 0.237342
R5125 VSS.n2759 VSS.n305 0.237342
R5126 VSS.n2760 VSS.n2759 0.237342
R5127 VSS.n2761 VSS.n2760 0.237342
R5128 VSS.n2761 VSS.n301 0.237342
R5129 VSS.n2767 VSS.n301 0.237342
R5130 VSS.n2768 VSS.n2767 0.237342
R5131 VSS.n2769 VSS.n2768 0.237342
R5132 VSS.n2769 VSS.n297 0.237342
R5133 VSS.n2775 VSS.n297 0.237342
R5134 VSS.n2776 VSS.n2775 0.237342
R5135 VSS.n2778 VSS.n2776 0.237342
R5136 VSS.n2778 VSS.n2777 0.237342
R5137 VSS.n2777 VSS.n293 0.237342
R5138 VSS.n2785 VSS.n293 0.237342
R5139 VSS.n2833 VSS.n2786 0.237342
R5140 VSS.n2827 VSS.n2786 0.237342
R5141 VSS.n2827 VSS.n2826 0.237342
R5142 VSS.n2826 VSS.n2825 0.237342
R5143 VSS.n2825 VSS.n2790 0.237342
R5144 VSS.n2819 VSS.n2790 0.237342
R5145 VSS.n2819 VSS.n2818 0.237342
R5146 VSS.n2818 VSS.n2817 0.237342
R5147 VSS.n2817 VSS.n2794 0.237342
R5148 VSS.n2811 VSS.n2794 0.237342
R5149 VSS.n2811 VSS.n2810 0.237342
R5150 VSS.n2810 VSS.n2809 0.237342
R5151 VSS.n2809 VSS.n2798 0.237342
R5152 VSS.n2803 VSS.n2798 0.237342
R5153 VSS.n2803 VSS.n2802 0.237342
R5154 VSS.n2802 VSS.n122 0.237342
R5155 VSS.n3098 VSS.n122 0.237342
R5156 VSS.n3098 VSS.n3097 0.237342
R5157 VSS.n3095 VSS.n125 0.237342
R5158 VSS.n3089 VSS.n125 0.237342
R5159 VSS.n3089 VSS.n3088 0.237342
R5160 VSS.n3088 VSS.n3087 0.237342
R5161 VSS.n3087 VSS.n132 0.237342
R5162 VSS.n134 VSS.n132 0.237342
R5163 VSS.n3080 VSS.n134 0.237342
R5164 VSS.n3080 VSS.n3079 0.237342
R5165 VSS.n3079 VSS.n3078 0.237342
R5166 VSS.n3078 VSS.n136 0.237342
R5167 VSS.n3072 VSS.n136 0.237342
R5168 VSS.n3072 VSS.n3071 0.237342
R5169 VSS.n3071 VSS.n3070 0.237342
R5170 VSS.n3070 VSS.n145 0.237342
R5171 VSS.n3064 VSS.n145 0.237342
R5172 VSS.n3064 VSS.n3063 0.237342
R5173 VSS.n3063 VSS.n3062 0.237342
R5174 VSS.n3062 VSS.n149 0.237342
R5175 VSS.n885 VSS.n884 0.237342
R5176 VSS.n884 VSS.n883 0.237342
R5177 VSS.n883 VSS.n833 0.237342
R5178 VSS.n877 VSS.n833 0.237342
R5179 VSS.n877 VSS.n876 0.237342
R5180 VSS.n876 VSS.n875 0.237342
R5181 VSS.n875 VSS.n836 0.237342
R5182 VSS.n869 VSS.n836 0.237342
R5183 VSS.n869 VSS.n868 0.237342
R5184 VSS.n868 VSS.n867 0.237342
R5185 VSS.n867 VSS.n841 0.237342
R5186 VSS.n861 VSS.n841 0.237342
R5187 VSS.n861 VSS.n860 0.237342
R5188 VSS.n860 VSS.n859 0.237342
R5189 VSS.n859 VSS.n843 0.237342
R5190 VSS.n854 VSS.n843 0.237342
R5191 VSS.n854 VSS.n853 0.237342
R5192 VSS.n853 VSS.n852 0.237342
R5193 VSS.n2170 VSS.n2169 0.237342
R5194 VSS.n2169 VSS.n2168 0.237342
R5195 VSS.n2168 VSS.n606 0.237342
R5196 VSS.n610 VSS.n606 0.237342
R5197 VSS.n2161 VSS.n610 0.237342
R5198 VSS.n2161 VSS.n2160 0.237342
R5199 VSS.n2160 VSS.n2159 0.237342
R5200 VSS.n2159 VSS.n611 0.237342
R5201 VSS.n1761 VSS.n611 0.237342
R5202 VSS.n2145 VSS.n1764 0.237342
R5203 VSS.n2145 VSS.n2144 0.237342
R5204 VSS.n2144 VSS.n2143 0.237342
R5205 VSS.n2143 VSS.n1765 0.237342
R5206 VSS.n2137 VSS.n1765 0.237342
R5207 VSS.n2137 VSS.n2136 0.237342
R5208 VSS.n2136 VSS.n2135 0.237342
R5209 VSS.n2135 VSS.n1769 0.237342
R5210 VSS.n2128 VSS.n2127 0.237342
R5211 VSS.n2127 VSS.n2126 0.237342
R5212 VSS.n2126 VSS.n1813 0.237342
R5213 VSS.n2120 VSS.n1813 0.237342
R5214 VSS.n2120 VSS.n2119 0.237342
R5215 VSS.n2119 VSS.n2118 0.237342
R5216 VSS.n2118 VSS.n1818 0.237342
R5217 VSS.n2112 VSS.n1818 0.237342
R5218 VSS.n2112 VSS.n2111 0.237342
R5219 VSS.n2111 VSS.n2110 0.237342
R5220 VSS.n2110 VSS.n1822 0.237342
R5221 VSS.n2104 VSS.n1822 0.237342
R5222 VSS.n2104 VSS.n2103 0.237342
R5223 VSS.n2103 VSS.n2102 0.237342
R5224 VSS.n2102 VSS.n1826 0.237342
R5225 VSS.n2096 VSS.n1826 0.237342
R5226 VSS.n2096 VSS.n2095 0.237342
R5227 VSS.n2095 VSS.n2094 0.237342
R5228 VSS.n1835 VSS.n1832 0.237342
R5229 VSS.n2046 VSS.n1835 0.237342
R5230 VSS.n2046 VSS.n2045 0.237342
R5231 VSS.n2045 VSS.n2044 0.237342
R5232 VSS.n2044 VSS.n1836 0.237342
R5233 VSS.n2038 VSS.n1836 0.237342
R5234 VSS.n2038 VSS.n2037 0.237342
R5235 VSS.n2037 VSS.n2036 0.237342
R5236 VSS.n2036 VSS.n1840 0.237342
R5237 VSS.n2030 VSS.n1840 0.237342
R5238 VSS.n2030 VSS.n2029 0.237342
R5239 VSS.n2029 VSS.n2028 0.237342
R5240 VSS.n2028 VSS.n1844 0.237342
R5241 VSS.n2022 VSS.n1844 0.237342
R5242 VSS.n2022 VSS.n2021 0.237342
R5243 VSS.n2021 VSS.n2020 0.237342
R5244 VSS.n2020 VSS.n1848 0.237342
R5245 VSS.n2014 VSS.n1848 0.237342
R5246 VSS.n2012 VSS.n1892 0.237342
R5247 VSS.n1896 VSS.n1892 0.237342
R5248 VSS.n2005 VSS.n1896 0.237342
R5249 VSS.n2005 VSS.n2004 0.237342
R5250 VSS.n2004 VSS.n2003 0.237342
R5251 VSS.n2003 VSS.n1897 0.237342
R5252 VSS.n1997 VSS.n1897 0.237342
R5253 VSS.n1997 VSS.n1996 0.237342
R5254 VSS.n1996 VSS.n1995 0.237342
R5255 VSS.n1995 VSS.n1901 0.237342
R5256 VSS.n1989 VSS.n1901 0.237342
R5257 VSS.n1989 VSS.n1988 0.237342
R5258 VSS.n1988 VSS.n1987 0.237342
R5259 VSS.n1987 VSS.n1905 0.237342
R5260 VSS.n1981 VSS.n1905 0.237342
R5261 VSS.n1981 VSS.n1980 0.237342
R5262 VSS.n1980 VSS.n1979 0.237342
R5263 VSS.n1979 VSS.n1909 0.237342
R5264 VSS.n1972 VSS.n1971 0.237342
R5265 VSS.n1971 VSS.n1970 0.237342
R5266 VSS.n1970 VSS.n1952 0.237342
R5267 VSS.n1964 VSS.n1952 0.237342
R5268 VSS.n1964 VSS.n1963 0.237342
R5269 VSS.n1963 VSS.n1962 0.237342
R5270 VSS.n1962 VSS.n1957 0.237342
R5271 VSS.n1957 VSS.n85 0.237342
R5272 VSS.n3155 VSS.n85 0.237342
R5273 VSS.n3155 VSS.n3154 0.237342
R5274 VSS.n3154 VSS.n3153 0.237342
R5275 VSS.n3153 VSS.n86 0.237342
R5276 VSS.n3147 VSS.n86 0.237342
R5277 VSS.n3147 VSS.n3146 0.237342
R5278 VSS.n3146 VSS.n3145 0.237342
R5279 VSS.n3145 VSS.n91 0.237342
R5280 VSS.n3139 VSS.n91 0.237342
R5281 VSS.n3139 VSS.n3138 0.237342
R5282 VSS.n3136 VSS.n96 0.237342
R5283 VSS.n3130 VSS.n96 0.237342
R5284 VSS.n3130 VSS.n3129 0.237342
R5285 VSS.n3129 VSS.n3128 0.237342
R5286 VSS.n3128 VSS.n102 0.237342
R5287 VSS.n3122 VSS.n102 0.237342
R5288 VSS.n3122 VSS.n3121 0.237342
R5289 VSS.n3121 VSS.n3120 0.237342
R5290 VSS.n3120 VSS.n106 0.237342
R5291 VSS.n3114 VSS.n106 0.237342
R5292 VSS.n3114 VSS.n3113 0.237342
R5293 VSS.n3113 VSS.n3112 0.237342
R5294 VSS.n3112 VSS.n109 0.237342
R5295 VSS.n3106 VSS.n109 0.237342
R5296 VSS.n3106 VSS.n3105 0.237342
R5297 VSS.n3105 VSS.n3104 0.237342
R5298 VSS.n3104 VSS.n114 0.237342
R5299 VSS.n745 VSS.n114 0.237342
R5300 VSS.n747 VSS.n698 0.237342
R5301 VSS.n753 VSS.n698 0.237342
R5302 VSS.n754 VSS.n753 0.237342
R5303 VSS.n755 VSS.n754 0.237342
R5304 VSS.n755 VSS.n696 0.237342
R5305 VSS.n696 VSS.n695 0.237342
R5306 VSS.n762 VSS.n695 0.237342
R5307 VSS.n763 VSS.n762 0.237342
R5308 VSS.n764 VSS.n763 0.237342
R5309 VSS.n764 VSS.n693 0.237342
R5310 VSS.n769 VSS.n693 0.237342
R5311 VSS.n770 VSS.n769 0.237342
R5312 VSS.n771 VSS.n770 0.237342
R5313 VSS.n771 VSS.n691 0.237342
R5314 VSS.n777 VSS.n691 0.237342
R5315 VSS.n778 VSS.n777 0.237342
R5316 VSS.n779 VSS.n778 0.237342
R5317 VSS.n779 VSS.n689 0.237342
R5318 VSS.n911 VSS.n910 0.237342
R5319 VSS.n912 VSS.n911 0.237342
R5320 VSS.n912 VSS.n686 0.237342
R5321 VSS.n918 VSS.n686 0.237342
R5322 VSS.n919 VSS.n918 0.237342
R5323 VSS.n920 VSS.n919 0.237342
R5324 VSS.n920 VSS.n684 0.237342
R5325 VSS.n926 VSS.n684 0.237342
R5326 VSS.n927 VSS.n926 0.237342
R5327 VSS.n928 VSS.n927 0.237342
R5328 VSS.n928 VSS.n682 0.237342
R5329 VSS.n934 VSS.n682 0.237342
R5330 VSS.n935 VSS.n934 0.237342
R5331 VSS.n936 VSS.n935 0.237342
R5332 VSS.n936 VSS.n680 0.237342
R5333 VSS.n942 VSS.n680 0.237342
R5334 VSS.n943 VSS.n942 0.237342
R5335 VSS.n944 VSS.n943 0.237342
R5336 VSS.n1553 VSS.n1552 0.237342
R5337 VSS.n1552 VSS.n1551 0.237342
R5338 VSS.n1551 VSS.n1449 0.237342
R5339 VSS.n1545 VSS.n1449 0.237342
R5340 VSS.n1545 VSS.n1544 0.237342
R5341 VSS.n1544 VSS.n1543 0.237342
R5342 VSS.n1543 VSS.n1509 0.237342
R5343 VSS.n1537 VSS.n1509 0.237342
R5344 VSS.n1535 VSS.n1534 0.237342
R5345 VSS.n1534 VSS.n1514 0.237342
R5346 VSS.n1528 VSS.n1514 0.237342
R5347 VSS.n1528 VSS.n1527 0.237342
R5348 VSS.n1527 VSS.n1526 0.237342
R5349 VSS.n1526 VSS.n1518 0.237342
R5350 VSS.n1520 VSS.n1518 0.237342
R5351 VSS.n1520 VSS.n531 0.237342
R5352 VSS.n2342 VSS.n531 0.237342
R5353 VSS.n2344 VSS.n526 0.237342
R5354 VSS.n2350 VSS.n526 0.237342
R5355 VSS.n2351 VSS.n2350 0.237342
R5356 VSS.n2352 VSS.n2351 0.237342
R5357 VSS.n2352 VSS.n522 0.237342
R5358 VSS.n2358 VSS.n522 0.237342
R5359 VSS.n2359 VSS.n2358 0.237342
R5360 VSS.n2362 VSS.n2359 0.237342
R5361 VSS.n2368 VSS.n518 0.237342
R5362 VSS.n2369 VSS.n2368 0.237342
R5363 VSS.n2370 VSS.n2369 0.237342
R5364 VSS.n2370 VSS.n514 0.237342
R5365 VSS.n2376 VSS.n514 0.237342
R5366 VSS.n2377 VSS.n2376 0.237342
R5367 VSS.n2378 VSS.n2377 0.237342
R5368 VSS.n2378 VSS.n510 0.237342
R5369 VSS.n2384 VSS.n510 0.237342
R5370 VSS.n2434 VSS.n2433 0.237342
R5371 VSS.n2433 VSS.n2432 0.237342
R5372 VSS.n2432 VSS.n2386 0.237342
R5373 VSS.n2426 VSS.n2386 0.237342
R5374 VSS.n2426 VSS.n2425 0.237342
R5375 VSS.n2425 VSS.n2424 0.237342
R5376 VSS.n2424 VSS.n2390 0.237342
R5377 VSS.n2418 VSS.n2390 0.237342
R5378 VSS.n2416 VSS.n2415 0.237342
R5379 VSS.n2415 VSS.n2395 0.237342
R5380 VSS.n2409 VSS.n2395 0.237342
R5381 VSS.n2409 VSS.n2408 0.237342
R5382 VSS.n2408 VSS.n2407 0.237342
R5383 VSS.n2407 VSS.n2399 0.237342
R5384 VSS.n2401 VSS.n2399 0.237342
R5385 VSS.n2401 VSS.n411 0.237342
R5386 VSS.n2609 VSS.n411 0.237342
R5387 VSS.n2611 VSS.n406 0.237342
R5388 VSS.n2617 VSS.n406 0.237342
R5389 VSS.n2618 VSS.n2617 0.237342
R5390 VSS.n2619 VSS.n2618 0.237342
R5391 VSS.n2619 VSS.n402 0.237342
R5392 VSS.n2625 VSS.n402 0.237342
R5393 VSS.n2626 VSS.n2625 0.237342
R5394 VSS.n2629 VSS.n2626 0.237342
R5395 VSS.n2635 VSS.n398 0.237342
R5396 VSS.n2636 VSS.n2635 0.237342
R5397 VSS.n2637 VSS.n2636 0.237342
R5398 VSS.n2637 VSS.n394 0.237342
R5399 VSS.n2643 VSS.n394 0.237342
R5400 VSS.n2644 VSS.n2643 0.237342
R5401 VSS.n2645 VSS.n2644 0.237342
R5402 VSS.n2645 VSS.n390 0.237342
R5403 VSS.n2651 VSS.n390 0.237342
R5404 VSS.n2706 VSS.n2705 0.237342
R5405 VSS.n2705 VSS.n2704 0.237342
R5406 VSS.n2704 VSS.n2653 0.237342
R5407 VSS.n2698 VSS.n2653 0.237342
R5408 VSS.n2698 VSS.n2697 0.237342
R5409 VSS.n2697 VSS.n2696 0.237342
R5410 VSS.n2696 VSS.n2657 0.237342
R5411 VSS.n2690 VSS.n2657 0.237342
R5412 VSS.n2688 VSS.n2687 0.237342
R5413 VSS.n2687 VSS.n2662 0.237342
R5414 VSS.n2681 VSS.n2662 0.237342
R5415 VSS.n2681 VSS.n2680 0.237342
R5416 VSS.n2680 VSS.n2679 0.237342
R5417 VSS.n2679 VSS.n2666 0.237342
R5418 VSS.n2673 VSS.n2666 0.237342
R5419 VSS.n2673 VSS.n2672 0.237342
R5420 VSS.n2672 VSS.n2671 0.237342
R5421 VSS.n2884 VSS.n2883 0.237342
R5422 VSS.n2885 VSS.n2884 0.237342
R5423 VSS.n2885 VSS.n260 0.237342
R5424 VSS.n2891 VSS.n260 0.237342
R5425 VSS.n2892 VSS.n2891 0.237342
R5426 VSS.n2893 VSS.n2892 0.237342
R5427 VSS.n2893 VSS.n256 0.237342
R5428 VSS.n2899 VSS.n256 0.237342
R5429 VSS.n2902 VSS.n2901 0.237342
R5430 VSS.n2902 VSS.n251 0.237342
R5431 VSS.n2908 VSS.n251 0.237342
R5432 VSS.n2909 VSS.n2908 0.237342
R5433 VSS.n2910 VSS.n2909 0.237342
R5434 VSS.n2910 VSS.n247 0.237342
R5435 VSS.n2916 VSS.n247 0.237342
R5436 VSS.n2917 VSS.n2916 0.237342
R5437 VSS.n2941 VSS.n2917 0.237342
R5438 VSS.n2939 VSS.n2926 0.237342
R5439 VSS.n2933 VSS.n2926 0.237342
R5440 VSS.n2933 VSS.n2932 0.237342
R5441 VSS.n2932 VSS.n2931 0.237342
R5442 VSS.n2931 VSS.n199 0.237342
R5443 VSS.n2965 VSS.n199 0.237342
R5444 VSS.n2966 VSS.n2965 0.237342
R5445 VSS.n2968 VSS.n2966 0.237342
R5446 VSS.n2968 VSS.n2967 0.237342
R5447 VSS.n2975 VSS.n2974 0.237342
R5448 VSS.n2976 VSS.n2975 0.237342
R5449 VSS.n2976 VSS.n190 0.237342
R5450 VSS.n2982 VSS.n190 0.237342
R5451 VSS.n2983 VSS.n2982 0.237342
R5452 VSS.n2984 VSS.n2983 0.237342
R5453 VSS.n2984 VSS.n186 0.237342
R5454 VSS.n2990 VSS.n186 0.237342
R5455 VSS.n3038 VSS.n3037 0.237342
R5456 VSS.n3037 VSS.n3036 0.237342
R5457 VSS.n3036 VSS.n2992 0.237342
R5458 VSS.n3030 VSS.n2992 0.237342
R5459 VSS.n3030 VSS.n3029 0.237342
R5460 VSS.n3029 VSS.n3028 0.237342
R5461 VSS.n3028 VSS.n2995 0.237342
R5462 VSS.n3022 VSS.n2995 0.237342
R5463 VSS.n3022 VSS.n3021 0.237342
R5464 VSS.n3021 VSS.n3020 0.237342
R5465 VSS.n3020 VSS.n3000 0.237342
R5466 VSS.n3014 VSS.n3000 0.237342
R5467 VSS.n3014 VSS.n3013 0.237342
R5468 VSS.n3013 VSS.n3012 0.237342
R5469 VSS.n3012 VSS.n3004 0.237342
R5470 VSS.n3006 VSS.n3004 0.237342
R5471 VSS.n3006 VSS.n2 0.237342
R5472 VSS.n3483 VSS.n2 0.237342
R5473 VSS.n2209 VSS.n596 0.235007
R5474 VSS.t190 VSS.n46 0.233316
R5475 VSS.n1693 VSS.n1692 0.229053
R5476 VSS.n1379 VSS.n1156 0.226684
R5477 VSS.n1641 VSS.n604 0.226498
R5478 VSS.n1147 VSS.n1146 0.223034
R5479 VSS.n1347 VSS.n1225 0.218395
R5480 VSS.n1261 VSS.n1260 0.218395
R5481 VSS.n3442 VSS.n3441 0.217142
R5482 VSS.n1373 VSS.n1204 0.207737
R5483 VSS.n1378 VSS.n1377 0.207737
R5484 VSS.n1579 VSS.n1578 0.207623
R5485 VSS.n1764 VSS.n1759 0.204184
R5486 VSS.n1650 VSS.n1079 0.1994
R5487 VSS.n1608 VSS.n1607 0.193093
R5488 VSS.n1607 VSS.n1606 0.193093
R5489 VSS.n33 VSS.n13 0.193093
R5490 VSS.n34 VSS.n33 0.193093
R5491 VSS.n3474 VSS.n3473 0.193093
R5492 VSS.n3475 VSS.n3474 0.193093
R5493 VSS.n1694 VSS.n1693 0.192342
R5494 VSS.n1057 VSS.n1056 0.189974
R5495 VSS.n1358 VSS.n1157 0.187417
R5496 VSS.n1246 VSS.n1216 0.186075
R5497 VSS.n1126 VSS.n1082 0.183582
R5498 VSS.n1438 VSS.n1414 0.183582
R5499 VSS.n1592 VSS.n1412 0.183582
R5500 VSS.n1116 VSS.n1110 0.183187
R5501 VSS.n2187 VSS.n597 0.181768
R5502 VSS.n1143 VSS.n1142 0.175877
R5503 VSS.n1386 VSS.n1151 0.1697
R5504 VSS.n1629 VSS.n1627 0.1661
R5505 VSS.n1632 VSS.n1631 0.1661
R5506 VSS.n41 VSS.n40 0.165427
R5507 VSS.n1433 VSS.n1432 0.163548
R5508 VSS.n3045 VSS.n3044 0.161553
R5509 VSS.n2299 VSS.n2252 0.161553
R5510 VSS.n2475 VSS.n2474 0.161553
R5511 VSS.n2566 VSS.n2514 0.161553
R5512 VSS.n361 VSS.n309 0.161553
R5513 VSS.n2834 VSS.n2833 0.161553
R5514 VSS.n3096 VSS.n3095 0.161553
R5515 VSS.n885 VSS.n832 0.161553
R5516 VSS.n1658 VSS.n1071 0.161553
R5517 VSS.n1497 VSS.n1448 0.161236
R5518 VSS.n1465 VSS.n594 0.156415
R5519 VSS.n1536 VSS.n1535 0.150895
R5520 VSS.n2361 VSS.n518 0.150895
R5521 VSS.n2417 VSS.n2416 0.150895
R5522 VSS.n2628 VSS.n398 0.150895
R5523 VSS.n2689 VSS.n2688 0.150895
R5524 VSS.n2901 VSS.n2900 0.150895
R5525 VSS.n1696 VSS.n630 0.148156
R5526 VSS.n2128 VSS.n1812 0.147342
R5527 VSS.n1832 VSS.n1830 0.147342
R5528 VSS.n2013 VSS.n2012 0.147342
R5529 VSS.n1972 VSS.n1951 0.147342
R5530 VSS.n3137 VSS.n3136 0.147342
R5531 VSS.n747 VSS.n746 0.147342
R5532 VSS.n910 VSS.n688 0.147342
R5533 VSS.n2344 VSS.n2343 0.147342
R5534 VSS.n2434 VSS.n2385 0.147342
R5535 VSS.n2611 VSS.n2610 0.147342
R5536 VSS.n2706 VSS.n2652 0.147342
R5537 VSS.n2883 VSS.n264 0.147342
R5538 VSS.n2940 VSS.n2939 0.147342
R5539 VSS.n3038 VSS.n2991 0.147342
R5540 VSS.n1214 VSS.n1204 0.144974
R5541 VSS.n1425 VSS.n1424 0.141048
R5542 VSS.n642 VSS.n620 0.14
R5543 VSS.n646 VSS.n642 0.14
R5544 VSS.n994 VSS.n646 0.14
R5545 VSS.n994 VSS.n993 0.14
R5546 VSS.n993 VSS.n992 0.14
R5547 VSS.n992 VSS.n647 0.14
R5548 VSS.n986 VSS.n647 0.14
R5549 VSS.n986 VSS.n985 0.14
R5550 VSS.n985 VSS.n984 0.14
R5551 VSS.n984 VSS.n653 0.14
R5552 VSS.n978 VSS.n653 0.14
R5553 VSS.n978 VSS.n977 0.14
R5554 VSS.n977 VSS.n976 0.14
R5555 VSS.n976 VSS.n671 0.14
R5556 VSS.n970 VSS.n671 0.14
R5557 VSS.n970 VSS.n969 0.14
R5558 VSS.n969 VSS.n968 0.14
R5559 VSS.n968 VSS.n949 0.14
R5560 VSS.n2974 VSS.n195 0.139053
R5561 VSS.n1437 VSS.n1436 0.13889
R5562 VSS.n1133 VSS.n1132 0.138582
R5563 VSS.n1429 VSS.n1428 0.138582
R5564 VSS.n1584 VSS.n1583 0.138582
R5565 VSS.n617 VSS.n616 0.137401
R5566 VSS.n1142 VSS.n1141 0.137349
R5567 VSS.n1215 VSS.n1214 0.13667
R5568 VSS.n1643 VSS.n1642 0.132545
R5569 VSS.n1379 VSS.n1378 0.131947
R5570 VSS.n1483 VSS.n593 0.128528
R5571 VSS.n1135 VSS.n1134 0.128411
R5572 VSS.n1812 VSS.n1769 0.128395
R5573 VSS.n2094 VSS.n1830 0.128395
R5574 VSS.n2014 VSS.n2013 0.128395
R5575 VSS.n1951 VSS.n1909 0.128395
R5576 VSS.n3138 VSS.n3137 0.128395
R5577 VSS.n746 VSS.n745 0.128395
R5578 VSS.n689 VSS.n688 0.128395
R5579 VSS.n2343 VSS.n2342 0.128395
R5580 VSS.n2385 VSS.n2384 0.128395
R5581 VSS.n2610 VSS.n2609 0.128395
R5582 VSS.n2652 VSS.n2651 0.128395
R5583 VSS.n2671 VSS.n264 0.128395
R5584 VSS.n2941 VSS.n2940 0.128395
R5585 VSS.n2991 VSS.n2990 0.128395
R5586 VSS.n1486 VSS.n593 0.125993
R5587 VSS.n1432 VSS.n1431 0.123479
R5588 VSS.n40 VSS.n27 0.120757
R5589 VSS.n1583 VSS.n1582 0.120089
R5590 VSS.n2211 VSS.n2210 0.118921
R5591 VSS.n1353 VSS.n1157 0.118667
R5592 VSS.n1427 VSS.n1426 0.117315
R5593 VSS.n1271 VSS.n1057 0.116553
R5594 VSS.n32 VSS.n26 0.114565
R5595 VSS.n1131 VSS.n1130 0.114233
R5596 VSS.n2252 VSS.n2251 0.114184
R5597 VSS.n2474 VSS.n2473 0.114184
R5598 VSS.n2514 VSS.n2513 0.114184
R5599 VSS.n2532 VSS.n361 0.114184
R5600 VSS.n2834 VSS.n2785 0.114184
R5601 VSS.n3097 VSS.n3096 0.114184
R5602 VSS.n832 VSS.n149 0.114184
R5603 VSS.n1580 VSS.n1579 0.113925
R5604 VSS.n678 VSS.n677 0.1085
R5605 VSS.n30 VSS.n29 0.108076
R5606 VSS.n3484 VSS.n0 0.106292
R5607 VSS.n1620 VSS.n1619 0.104969
R5608 VSS.n2170 VSS.n595 0.104711
R5609 VSS.n1553 VSS.n1448 0.104711
R5610 VSS.n1435 VSS.n1434 0.10437
R5611 VSS.n2940 VSS.n2925 0.102342
R5612 VSS.n2991 VSS.n185 0.102342
R5613 VSS.n2343 VSS.n530 0.102342
R5614 VSS.n2385 VSS.n509 0.102342
R5615 VSS.n2610 VSS.n410 0.102342
R5616 VSS.n2652 VSS.n389 0.102342
R5617 VSS.n2872 VSS.n264 0.102342
R5618 VSS.n3096 VSS.n123 0.101158
R5619 VSS.n2252 VSS.n567 0.101158
R5620 VSS.n2474 VSS.n468 0.101158
R5621 VSS.n2514 VSS.n446 0.101158
R5622 VSS.n2742 VSS.n361 0.101158
R5623 VSS.n2838 VSS.n2834 0.101158
R5624 VSS.n832 VSS.n831 0.101158
R5625 VSS.n2967 VSS.n195 0.0987895
R5626 VSS.n2194 VSS.n594 0.0981056
R5627 VSS.n1618 VSS.n1617 0.0971559
R5628 VSS.n1264 VSS.n1225 0.0952368
R5629 VSS.n1308 VSS.n1261 0.0952368
R5630 VSS.n3464 VSS.n3463 0.095011
R5631 VSS.n1354 VSS.n1353 0.0948615
R5632 VSS.n1570 VSS.n1569 0.0941986
R5633 VSS.n1107 VSS.n1106 0.0933571
R5634 VSS.n1605 VSS.n1107 0.0933571
R5635 VSS.n1611 VSS.n1610 0.0933571
R5636 VSS.n1612 VSS.n1611 0.0933571
R5637 VSS.n1614 VSS.n1613 0.0933571
R5638 VSS.n1613 VSS.n1612 0.0933571
R5639 VSS.n1391 VSS.n1149 0.0933571
R5640 VSS.n1391 VSS.n1390 0.0933571
R5641 VSS.n3450 VSS.n3449 0.0933571
R5642 VSS.n3451 VSS.n3450 0.0933571
R5643 VSS.n3458 VSS.n3457 0.0933571
R5644 VSS.n3459 VSS.n3458 0.0933571
R5645 VSS.n3461 VSS.n3460 0.0933571
R5646 VSS.n3460 VSS.n3459 0.0933571
R5647 VSS.n3470 VSS.n3469 0.0933571
R5648 VSS.n3469 VSS.n3468 0.0933571
R5649 VSS.n3479 VSS.n0 0.0933571
R5650 VSS.n3480 VSS.n3479 0.0933571
R5651 VSS.n1424 VSS.n1422 0.0905
R5652 VSS.n322 VSS.n68 0.0895206
R5653 VSS.n3442 VSS.n43 0.0874537
R5654 VSS.n2153 VSS.n618 0.0874227
R5655 VSS.n1537 VSS.n1536 0.0869474
R5656 VSS.n2362 VSS.n2361 0.0869474
R5657 VSS.n2418 VSS.n2417 0.0869474
R5658 VSS.n2629 VSS.n2628 0.0869474
R5659 VSS.n2690 VSS.n2689 0.0869474
R5660 VSS.n2900 VSS.n2899 0.0869474
R5661 VSS.n746 VSS.n742 0.0833947
R5662 VSS.n3137 VSS.n95 0.0833947
R5663 VSS.n1951 VSS.n1950 0.0833947
R5664 VSS.n2013 VSS.n1891 0.0833947
R5665 VSS.n1812 VSS.n1811 0.0833947
R5666 VSS.n2057 VSS.n1830 0.0833947
R5667 VSS.n784 VSS.n688 0.0833947
R5668 VSS.n1567 VSS.n1566 0.0831718
R5669 VSS.n1395 VSS.n1394 0.0821077
R5670 VSS.n1694 VSS.n1056 0.08159
R5671 VSS.n1129 VSS.n1128 0.0797123
R5672 VSS.n1353 VSS.n1150 0.0772371
R5673 VSS.n1117 VSS.n1109 0.0755346
R5674 VSS.n1636 VSS.n1632 0.0743
R5675 VSS.n1636 VSS.n1635 0.0743
R5676 VSS.n1646 VSS.n1080 0.0743
R5677 VSS.n1647 VSS.n1646 0.0743
R5678 VSS.n2208 VSS.n597 0.0727535
R5679 VSS.n1400 VSS.n1396 0.0711109
R5680 VSS.n1146 VSS.n1145 0.0695411
R5681 VSS.n1436 VSS.n1435 0.0692329
R5682 VSS.n1649 VSS.n1648 0.0689
R5683 VSS.n1359 VSS.n1358 0.0680325
R5684 VSS.n1360 VSS.n1359 0.0680325
R5685 VSS.n1113 VSS.n1083 0.0680325
R5686 VSS.n1638 VSS.n1083 0.0680325
R5687 VSS.n1396 VSS.n1395 0.0653232
R5688 VSS.n1399 VSS.n1398 0.0653232
R5689 VSS.n1398 VSS.n1101 0.0653232
R5690 VSS.n1616 VSS.n1615 0.0653232
R5691 VSS.n1619 VSS.n1618 0.0653232
R5692 VSS.n27 VSS.n22 0.0626638
R5693 VSS.n1755 VSS.n636 0.0626562
R5694 VSS.n1431 VSS.n1430 0.060911
R5695 VSS.n1128 VSS.n1127 0.0596781
R5696 VSS.n1422 VSS.n1421 0.0596781
R5697 VSS.n1130 VSS.n1129 0.0593699
R5698 VSS.n1144 VSS.n1143 0.0584452
R5699 VSS.n1140 VSS.n1139 0.0584452
R5700 VSS.n1137 VSS.n1136 0.0584452
R5701 VSS.n1127 VSS.n1126 0.0584452
R5702 VSS.n1430 VSS.n1429 0.0584452
R5703 VSS.n1438 VSS.n1437 0.0584452
R5704 VSS.n1578 VSS.n1412 0.0584452
R5705 VSS.n3484 VSS.n1 0.0576584
R5706 VSS.n2154 VSS.n615 0.0561818
R5707 VSS.n1139 VSS.n1138 0.0559795
R5708 VSS.n1136 VSS.n1135 0.0559795
R5709 VSS.n1571 VSS.n1570 0.0559795
R5710 VSS.n1595 VSS.n1594 0.0559198
R5711 VSS.n1615 VSS.n1614 0.05259
R5712 VSS.n3447 VSS.n28 0.0519837
R5713 VSS.n1566 VSS.n1565 0.0517977
R5714 VSS.n1565 VSS.n1564 0.0517977
R5715 VSS.n1564 VSS.n1563 0.0517977
R5716 VSS.n1563 VSS.n1408 0.0517977
R5717 VSS.n1599 VSS.n1598 0.0517977
R5718 VSS.n1597 VSS.n1596 0.0517977
R5719 VSS.n1596 VSS.n1595 0.0517977
R5720 VSS.n1600 VSS.n1408 0.0513397
R5721 VSS.n1693 VSS.n1057 0.0490526
R5722 VSS.n2151 VSS.n2150 0.0480786
R5723 VSS.n1115 VSS.n1114 0.0470589
R5724 VSS.n1112 VSS.n1111 0.0470589
R5725 VSS.n1087 VSS.n1086 0.0470589
R5726 VSS.n1086 VSS.n1085 0.0470589
R5727 VSS.n1085 VSS.n1084 0.0470589
R5728 VSS.n1084 VSS.n1081 0.0470589
R5729 VSS.n3096 VSS.n124 0.0466842
R5730 VSS.n2834 VSS.n292 0.0466842
R5731 VSS.n1922 VSS.n361 0.0466842
R5732 VSS.n2514 VSS.n447 0.0466842
R5733 VSS.n2252 VSS.n568 0.0466842
R5734 VSS.n2474 VSS.n469 0.0466842
R5735 VSS.n832 VSS.n813 0.0466842
R5736 VSS.n3445 VSS.n3444 0.0461627
R5737 VSS.n1116 VSS.n1115 0.0459157
R5738 VSS.n1114 VSS.n1113 0.0438372
R5739 VSS.n1640 VSS.n1088 0.0438333
R5740 VSS.n1640 VSS.n1639 0.0438333
R5741 VSS.n1601 VSS.n1600 0.0438333
R5742 VSS.n1602 VSS.n1601 0.0438333
R5743 VSS.n1696 VSS.n1695 0.0423279
R5744 VSS.n1620 VSS.n1095 0.03875
R5745 VSS.n1400 VSS.n1399 0.0386994
R5746 VSS.n1755 VSS.n635 0.035375
R5747 VSS.n998 VSS.n636 0.035375
R5748 VSS.n998 VSS.n997 0.035375
R5749 VSS.n997 VSS.n996 0.035375
R5750 VSS.n996 VSS.n643 0.035375
R5751 VSS.n990 VSS.n643 0.035375
R5752 VSS.n990 VSS.n989 0.035375
R5753 VSS.n989 VSS.n988 0.035375
R5754 VSS.n988 VSS.n650 0.035375
R5755 VSS.n982 VSS.n650 0.035375
R5756 VSS.n982 VSS.n981 0.035375
R5757 VSS.n981 VSS.n980 0.035375
R5758 VSS.n980 VSS.n668 0.035375
R5759 VSS.n974 VSS.n668 0.035375
R5760 VSS.n974 VSS.n973 0.035375
R5761 VSS.n973 VSS.n972 0.035375
R5762 VSS.n972 VSS.n674 0.035375
R5763 VSS.n1761 VSS.n1759 0.0336579
R5764 VSS.n1568 VSS.n1096 0.032
R5765 VSS.n3440 VSS.t190 0.0317616
R5766 VSS.n3464 VSS.n3462 0.0317469
R5767 VSS.n1621 VSS.n1620 0.0314524
R5768 VSS.n1622 VSS.n1621 0.0314524
R5769 VSS.n1591 VSS.n1590 0.0314524
R5770 VSS.n1590 VSS.n1589 0.0314524
R5771 VSS.n3274 VSS.n3237 0.0303125
R5772 VSS.n3270 VSS.n3237 0.0303125
R5773 VSS.n3270 VSS.n3269 0.0303125
R5774 VSS.n3269 VSS.n3268 0.0303125
R5775 VSS.n3268 VSS.n3239 0.0303125
R5776 VSS.n3264 VSS.n3239 0.0303125
R5777 VSS.n3264 VSS.n3263 0.0303125
R5778 VSS.n3263 VSS.n3262 0.0303125
R5779 VSS.n3262 VSS.n3241 0.0303125
R5780 VSS.n3258 VSS.n3241 0.0303125
R5781 VSS.n3258 VSS.n3257 0.0303125
R5782 VSS.n3257 VSS.n3256 0.0303125
R5783 VSS.n3256 VSS.n3243 0.0303125
R5784 VSS.n3252 VSS.n3243 0.0303125
R5785 VSS.n3252 VSS.n3251 0.0303125
R5786 VSS.n3251 VSS.n3250 0.0303125
R5787 VSS.n3250 VSS.n3245 0.0303125
R5788 VSS.n3246 VSS.n3245 0.0303125
R5789 VSS.n3246 VSS.n43 0.0303125
R5790 VSS.n3273 VSS.n3272 0.0303125
R5791 VSS.n3272 VSS.n3271 0.0303125
R5792 VSS.n3271 VSS.n3238 0.0303125
R5793 VSS.n3267 VSS.n3238 0.0303125
R5794 VSS.n3267 VSS.n3266 0.0303125
R5795 VSS.n3266 VSS.n3265 0.0303125
R5796 VSS.n3265 VSS.n3240 0.0303125
R5797 VSS.n3261 VSS.n3240 0.0303125
R5798 VSS.n3261 VSS.n3260 0.0303125
R5799 VSS.n3260 VSS.n3259 0.0303125
R5800 VSS.n3259 VSS.n3242 0.0303125
R5801 VSS.n3255 VSS.n3242 0.0303125
R5802 VSS.n3255 VSS.n3254 0.0303125
R5803 VSS.n3254 VSS.n3253 0.0303125
R5804 VSS.n3253 VSS.n3244 0.0303125
R5805 VSS.n3249 VSS.n3244 0.0303125
R5806 VSS.n3249 VSS.n3248 0.0303125
R5807 VSS.n3248 VSS.n3247 0.0303125
R5808 VSS.n3247 VSS.n44 0.0303125
R5809 VSS.n3441 VSS.n44 0.0303125
R5810 VSS.n1428 VSS.n1427 0.030089
R5811 VSS.n1354 VSS.n1089 0.0300285
R5812 VSS.n3441 VSS.n3440 0.0299118
R5813 VSS.n3044 VSS.n162 0.0289211
R5814 VSS.n1117 VSS.n1116 0.028664
R5815 VSS.n1001 VSS.n640 0.0284
R5816 VSS.n655 VSS.n640 0.0284
R5817 VSS.n655 VSS.n644 0.0284
R5818 VSS.n658 VSS.n644 0.0284
R5819 VSS.n658 VSS.n648 0.0284
R5820 VSS.n661 VSS.n648 0.0284
R5821 VSS.n661 VSS.n651 0.0284
R5822 VSS.n665 VSS.n651 0.0284
R5823 VSS.n666 VSS.n665 0.0284
R5824 VSS.n951 VSS.n666 0.0284
R5825 VSS.n951 VSS.n669 0.0284
R5826 VSS.n954 VSS.n669 0.0284
R5827 VSS.n954 VSS.n672 0.0284
R5828 VSS.n957 VSS.n672 0.0284
R5829 VSS.n957 VSS.n675 0.0284
R5830 VSS.n960 VSS.n675 0.0284
R5831 VSS.n960 VSS.n950 0.0284
R5832 VSS.n964 VSS.n950 0.0284
R5833 VSS.n1000 VSS.n999 0.0284
R5834 VSS.n999 VSS.n641 0.0284
R5835 VSS.n995 VSS.n641 0.0284
R5836 VSS.n995 VSS.n645 0.0284
R5837 VSS.n991 VSS.n645 0.0284
R5838 VSS.n991 VSS.n649 0.0284
R5839 VSS.n987 VSS.n649 0.0284
R5840 VSS.n987 VSS.n652 0.0284
R5841 VSS.n983 VSS.n652 0.0284
R5842 VSS.n983 VSS.n667 0.0284
R5843 VSS.n979 VSS.n667 0.0284
R5844 VSS.n979 VSS.n670 0.0284
R5845 VSS.n975 VSS.n670 0.0284
R5846 VSS.n975 VSS.n673 0.0284
R5847 VSS.n971 VSS.n673 0.0284
R5848 VSS.n971 VSS.n676 0.0284
R5849 VSS.n967 VSS.n676 0.0284
R5850 VSS.n1088 VSS.n1087 0.0279365
R5851 VSS.n3279 VSS.n3278 0.0274686
R5852 VSS.n1617 VSS.n1616 0.0271238
R5853 VSS.n1212 VSS.n1150 0.02642
R5854 VSS.n1364 VSS.n1215 0.0258274
R5855 VSS.n1138 VSS.n1137 0.0251575
R5856 VSS.n1132 VSS.n1131 0.0248493
R5857 VSS.n3477 VSS.n8 0.0245741
R5858 VSS.n3477 VSS.n3476 0.0245741
R5859 VSS.n1001 VSS.n639 0.0239
R5860 VSS.n1000 VSS.n628 0.0239
R5861 VSS.n1414 VSS.n1413 0.023
R5862 VSS.n3443 VSS.n3442 0.0229864
R5863 VSS.n1598 VSS.n1597 0.0220267
R5864 VSS.n1594 VSS.n1593 0.0220267
R5865 VSS.n656 VSS.n654 0.0219615
R5866 VSS.n657 VSS.n656 0.0219615
R5867 VSS.n659 VSS.n657 0.0219615
R5868 VSS.n660 VSS.n659 0.0219615
R5869 VSS.n662 VSS.n660 0.0219615
R5870 VSS.n663 VSS.n662 0.0219615
R5871 VSS.n664 VSS.n663 0.0219615
R5872 VSS.n664 VSS.t338 0.0219615
R5873 VSS.n952 VSS.t338 0.0219615
R5874 VSS.n953 VSS.n952 0.0219615
R5875 VSS.n955 VSS.n953 0.0219615
R5876 VSS.n956 VSS.n955 0.0219615
R5877 VSS.n958 VSS.n956 0.0219615
R5878 VSS.n959 VSS.n958 0.0219615
R5879 VSS.n961 VSS.n959 0.0219615
R5880 VSS.n962 VSS.n961 0.0219615
R5881 VSS.n963 VSS.n962 0.0219615
R5882 VSS.n1758 VSS.n621 0.0215938
R5883 VSS.n1643 VSS.n1081 0.0200381
R5884 VSS.n3434 VSS.n66 0.0199425
R5885 VSS.n3406 VSS.n66 0.0199425
R5886 VSS.n3413 VSS.n3406 0.0199425
R5887 VSS.n3414 VSS.n3413 0.0199425
R5888 VSS.n3415 VSS.n3414 0.0199425
R5889 VSS.n3415 VSS.n3403 0.0199425
R5890 VSS.n3421 VSS.n3403 0.0199425
R5891 VSS.n3421 VSS.n3170 0.0199425
R5892 VSS.n3425 VSS.n3170 0.0199425
R5893 VSS.n3425 VSS.n3401 0.0199425
R5894 VSS.n3401 VSS.n3400 0.0199425
R5895 VSS.n3400 VSS.n3171 0.0199425
R5896 VSS.n3175 VSS.n3171 0.0199425
R5897 VSS.n3392 VSS.n3175 0.0199425
R5898 VSS.n3392 VSS.n3176 0.0199425
R5899 VSS.n3388 VSS.n3176 0.0199425
R5900 VSS.n3388 VSS.n3179 0.0199425
R5901 VSS.n3382 VSS.n3179 0.0199425
R5902 VSS.n3382 VSS.n3381 0.0199425
R5903 VSS.n3381 VSS.n3183 0.0199425
R5904 VSS.n3377 VSS.n3183 0.0199425
R5905 VSS.n3377 VSS.n3185 0.0199425
R5906 VSS.n3188 VSS.n3185 0.0199425
R5907 VSS.n3191 VSS.n3188 0.0199425
R5908 VSS.n3366 VSS.n3191 0.0199425
R5909 VSS.n3366 VSS.n3192 0.0199425
R5910 VSS.n3362 VSS.n3192 0.0199425
R5911 VSS.n3362 VSS.n3194 0.0199425
R5912 VSS.n3356 VSS.n3194 0.0199425
R5913 VSS.n3356 VSS.n3354 0.0199425
R5914 VSS.n3354 VSS.n3353 0.0199425
R5915 VSS.n3353 VSS.n3197 0.0199425
R5916 VSS.n3347 VSS.n3197 0.0199425
R5917 VSS.n3347 VSS.n3201 0.0199425
R5918 VSS.n3343 VSS.n3201 0.0199425
R5919 VSS.n3343 VSS.n3204 0.0199425
R5920 VSS.n3206 VSS.n3204 0.0199425
R5921 VSS.n3209 VSS.n3206 0.0199425
R5922 VSS.n3332 VSS.n3209 0.0199425
R5923 VSS.n3332 VSS.n3210 0.0199425
R5924 VSS.n3328 VSS.n3210 0.0199425
R5925 VSS.n3328 VSS.n3212 0.0199425
R5926 VSS.n3322 VSS.n3212 0.0199425
R5927 VSS.n3322 VSS.n3321 0.0199425
R5928 VSS.n3321 VSS.n3320 0.0199425
R5929 VSS.n3320 VSS.n3215 0.0199425
R5930 VSS.n3314 VSS.n3215 0.0199425
R5931 VSS.n3314 VSS.n3220 0.0199425
R5932 VSS.n3310 VSS.n3220 0.0199425
R5933 VSS.n3310 VSS.n3222 0.0199425
R5934 VSS.n3224 VSS.n3222 0.0199425
R5935 VSS.n3227 VSS.n3224 0.0199425
R5936 VSS.n3299 VSS.n3227 0.0199425
R5937 VSS.n3299 VSS.n3228 0.0199425
R5938 VSS.n3295 VSS.n3228 0.0199425
R5939 VSS.n3295 VSS.n3230 0.0199425
R5940 VSS.n3289 VSS.n3230 0.0199425
R5941 VSS.n3289 VSS.n3288 0.0199425
R5942 VSS.n3288 VSS.n3234 0.0199425
R5943 VSS.n3284 VSS.n3234 0.0199425
R5944 VSS.n3284 VSS.n45 0.0199425
R5945 VSS.n3433 VSS.n67 0.0199425
R5946 VSS.n3409 VSS.n67 0.0199425
R5947 VSS.n3412 VSS.n3409 0.0199425
R5948 VSS.n3412 VSS.n3405 0.0199425
R5949 VSS.n3416 VSS.n3405 0.0199425
R5950 VSS.n3416 VSS.n3404 0.0199425
R5951 VSS.n3420 VSS.n3404 0.0199425
R5952 VSS.n3420 VSS.n3168 0.0199425
R5953 VSS.n3426 VSS.n3168 0.0199425
R5954 VSS.n3426 VSS.n3169 0.0199425
R5955 VSS.n3399 VSS.n3169 0.0199425
R5956 VSS.n3399 VSS.n3397 0.0199425
R5957 VSS.n3397 VSS.n3172 0.0199425
R5958 VSS.n3393 VSS.n3172 0.0199425
R5959 VSS.n3393 VSS.n3174 0.0199425
R5960 VSS.n3387 VSS.n3174 0.0199425
R5961 VSS.n3387 VSS.n3180 0.0199425
R5962 VSS.n3383 VSS.n3180 0.0199425
R5963 VSS.n3383 VSS.n3182 0.0199425
R5964 VSS.n3186 VSS.n3182 0.0199425
R5965 VSS.n3376 VSS.n3186 0.0199425
R5966 VSS.n3376 VSS.n3372 0.0199425
R5967 VSS.n3372 VSS.n3371 0.0199425
R5968 VSS.n3371 VSS.n3187 0.0199425
R5969 VSS.n3367 VSS.n3187 0.0199425
R5970 VSS.n3367 VSS.n3190 0.0199425
R5971 VSS.n3361 VSS.n3190 0.0199425
R5972 VSS.n3361 VSS.n3195 0.0199425
R5973 VSS.n3357 VSS.n3195 0.0199425
R5974 VSS.n3357 VSS.n3196 0.0199425
R5975 VSS.n3352 VSS.n3196 0.0199425
R5976 VSS.n3352 VSS.n3198 0.0199425
R5977 VSS.n3348 VSS.n3198 0.0199425
R5978 VSS.n3348 VSS.n3200 0.0199425
R5979 VSS.n3342 VSS.n3200 0.0199425
R5980 VSS.n3342 VSS.n3338 0.0199425
R5981 VSS.n3338 VSS.n3337 0.0199425
R5982 VSS.n3337 VSS.n3205 0.0199425
R5983 VSS.n3333 VSS.n3205 0.0199425
R5984 VSS.n3333 VSS.n3208 0.0199425
R5985 VSS.n3327 VSS.n3208 0.0199425
R5986 VSS.n3327 VSS.n3213 0.0199425
R5987 VSS.n3323 VSS.n3213 0.0199425
R5988 VSS.n3323 VSS.n3214 0.0199425
R5989 VSS.n3319 VSS.n3214 0.0199425
R5990 VSS.n3319 VSS.n3217 0.0199425
R5991 VSS.n3315 VSS.n3217 0.0199425
R5992 VSS.n3315 VSS.n3219 0.0199425
R5993 VSS.n3309 VSS.n3219 0.0199425
R5994 VSS.n3309 VSS.n3305 0.0199425
R5995 VSS.n3305 VSS.n3304 0.0199425
R5996 VSS.n3304 VSS.n3223 0.0199425
R5997 VSS.n3300 VSS.n3223 0.0199425
R5998 VSS.n3300 VSS.n3226 0.0199425
R5999 VSS.n3294 VSS.n3226 0.0199425
R6000 VSS.n3294 VSS.n3231 0.0199425
R6001 VSS.n3290 VSS.n3231 0.0199425
R6002 VSS.n3290 VSS.n3233 0.0199425
R6003 VSS.n3235 VSS.n3233 0.0199425
R6004 VSS.n3283 VSS.n3235 0.0199425
R6005 VSS.n3283 VSS.n3279 0.0199425
R6006 VSS.n1697 VSS.n1696 0.0198648
R6007 VSS.n1111 VSS.n1088 0.0196224
R6008 VSS.n2209 VSS.n2208 0.0195141
R6009 VSS.n654 VSS.t338 0.0191923
R6010 VSS.n1695 VSS.n1055 0.0189426
R6011 VSS.n948 VSS.n947 0.0188746
R6012 VSS.n947 VSS.n82 0.0188746
R6013 VSS.n629 VSS.n626 0.0183702
R6014 VSS.n638 VSS.n626 0.0183702
R6015 VSS.n631 VSS.n625 0.0183702
R6016 VSS.n637 VSS.n625 0.0183702
R6017 VSS.n633 VSS.n621 0.0183702
R6018 VSS.n1757 VSS.n623 0.0183702
R6019 VSS.n638 VSS.n632 0.0183702
R6020 VSS.n637 VSS.n634 0.0183702
R6021 VSS.n635 VSS.n623 0.0183702
R6022 VSS.n630 VSS.n629 0.0183702
R6023 VSS.n632 VSS.n631 0.0183702
R6024 VSS.n634 VSS.n633 0.0183702
R6025 VSS.n3275 VSS.n42 0.0183274
R6026 VSS.n3432 VSS.n3431 0.0176692
R6027 VSS.n3411 VSS.n69 0.0176692
R6028 VSS.n3411 VSS.n3410 0.0176692
R6029 VSS.n3418 VSS.n3417 0.0176692
R6030 VSS.n3419 VSS.n3418 0.0176692
R6031 VSS.n3419 VSS.n3166 0.0176692
R6032 VSS.n3427 VSS.n3167 0.0176692
R6033 VSS.n3398 VSS.n3167 0.0176692
R6034 VSS.n3396 VSS.n3395 0.0176692
R6035 VSS.n3395 VSS.n3394 0.0176692
R6036 VSS.n3394 VSS.n3173 0.0176692
R6037 VSS.n3386 VSS.n3385 0.0176692
R6038 VSS.n3385 VSS.n3384 0.0176692
R6039 VSS.n3384 VSS.n3181 0.0176692
R6040 VSS.n3373 VSS.n3181 0.0176692
R6041 VSS.n3375 VSS.n3373 0.0176692
R6042 VSS.n3375 VSS.n3374 0.0176692
R6043 VSS.n3370 VSS.n3369 0.0176692
R6044 VSS.n3369 VSS.n3368 0.0176692
R6045 VSS.n3368 VSS.n3189 0.0176692
R6046 VSS.n3360 VSS.n3359 0.0176692
R6047 VSS.n3359 VSS.n3358 0.0176692
R6048 VSS.n3351 VSS.n3199 0.0176692
R6049 VSS.n3351 VSS.n3350 0.0176692
R6050 VSS.n3350 VSS.n3349 0.0176692
R6051 VSS.n3341 VSS.n3339 0.0176692
R6052 VSS.n3341 VSS.n3340 0.0176692
R6053 VSS.n3336 VSS.n3335 0.0176692
R6054 VSS.n3335 VSS.n3334 0.0176692
R6055 VSS.n3334 VSS.n3207 0.0176692
R6056 VSS.n3326 VSS.n3325 0.0176692
R6057 VSS.n3325 VSS.n3324 0.0176692
R6058 VSS.n3318 VSS.n3218 0.0176692
R6059 VSS.n3318 VSS.n3317 0.0176692
R6060 VSS.n3317 VSS.n3316 0.0176692
R6061 VSS.n3308 VSS.n3306 0.0176692
R6062 VSS.n3308 VSS.n3307 0.0176692
R6063 VSS.n3303 VSS.n3302 0.0176692
R6064 VSS.n3302 VSS.n3301 0.0176692
R6065 VSS.n3301 VSS.n3225 0.0176692
R6066 VSS.n3293 VSS.n3292 0.0176692
R6067 VSS.n3292 VSS.n3291 0.0176692
R6068 VSS.n3291 VSS.n3232 0.0176692
R6069 VSS.n3282 VSS.n3280 0.0176692
R6070 VSS.n3282 VSS.n3281 0.0176692
R6071 VSS.n3307 VSS.n77 0.0173923
R6072 VSS.n3278 VSS.n3236 0.0171202
R6073 VSS.n3398 VSS.n72 0.0168385
R6074 VSS.n3435 VSS.n65 0.0165807
R6075 VSS.n3407 VSS.n65 0.0165807
R6076 VSS.n3408 VSS.n3407 0.0165807
R6077 VSS.n3408 VSS.n63 0.0165807
R6078 VSS.n3402 VSS.n64 0.0165807
R6079 VSS.n3422 VSS.n3402 0.0165807
R6080 VSS.n3423 VSS.n3422 0.0165807
R6081 VSS.n3424 VSS.n3423 0.0165807
R6082 VSS.n3424 VSS.n61 0.0165807
R6083 VSS.n3177 VSS.n62 0.0165807
R6084 VSS.n3178 VSS.n3177 0.0165807
R6085 VSS.n3391 VSS.n3178 0.0165807
R6086 VSS.n3391 VSS.n3390 0.0165807
R6087 VSS.n3390 VSS.n3389 0.0165807
R6088 VSS.n3389 VSS.n59 0.0165807
R6089 VSS.n3380 VSS.n60 0.0165807
R6090 VSS.n3380 VSS.n3379 0.0165807
R6091 VSS.n3379 VSS.n3378 0.0165807
R6092 VSS.n3378 VSS.n3184 0.0165807
R6093 VSS.n3184 VSS.n57 0.0165807
R6094 VSS.n3365 VSS.n58 0.0165807
R6095 VSS.n3365 VSS.n3364 0.0165807
R6096 VSS.n3364 VSS.n3363 0.0165807
R6097 VSS.n3363 VSS.n3193 0.0165807
R6098 VSS.n3355 VSS.n3193 0.0165807
R6099 VSS.n3355 VSS.n55 0.0165807
R6100 VSS.n3202 VSS.n56 0.0165807
R6101 VSS.n3346 VSS.n3202 0.0165807
R6102 VSS.n3346 VSS.n3345 0.0165807
R6103 VSS.n3345 VSS.n3344 0.0165807
R6104 VSS.n3344 VSS.n3203 0.0165807
R6105 VSS.n3203 VSS.n53 0.0165807
R6106 VSS.n3331 VSS.n54 0.0165807
R6107 VSS.n3331 VSS.n3330 0.0165807
R6108 VSS.n3330 VSS.n3329 0.0165807
R6109 VSS.n3329 VSS.n3211 0.0165807
R6110 VSS.n3211 VSS.n51 0.0165807
R6111 VSS.n3216 VSS.n52 0.0165807
R6112 VSS.n3221 VSS.n3216 0.0165807
R6113 VSS.n3313 VSS.n3221 0.0165807
R6114 VSS.n3313 VSS.n3312 0.0165807
R6115 VSS.n3312 VSS.n3311 0.0165807
R6116 VSS.n3311 VSS.n49 0.0165807
R6117 VSS.n3229 VSS.n50 0.0165807
R6118 VSS.n3298 VSS.n3229 0.0165807
R6119 VSS.n3298 VSS.n3297 0.0165807
R6120 VSS.n3297 VSS.n3296 0.0165807
R6121 VSS.n3296 VSS.n47 0.0165807
R6122 VSS.n3287 VSS.n48 0.0165807
R6123 VSS.n3287 VSS.n3286 0.0165807
R6124 VSS.n3286 VSS.n3285 0.0165807
R6125 VSS.n3285 VSS.n46 0.0165807
R6126 VSS.n3280 VSS.n78 0.0162846
R6127 VSS.n2154 VSS.n2153 0.0159762
R6128 VSS.n2155 VSS.n2154 0.0159762
R6129 VSS.t189 VSS.n64 0.0158026
R6130 VSS.t190 VSS.n47 0.0158026
R6131 VSS.n3324 VSS.n76 0.0157308
R6132 VSS.n3472 VSS.n8 0.0154357
R6133 VSS.n3410 VSS.n71 0.0151769
R6134 VSS.n3360 VSS.n3164 0.0151769
R6135 VSS.n3277 VSS.n3276 0.0151769
R6136 VSS.n3462 VSS.n22 0.0151333
R6137 VSS.n966 VSS.n965 0.0149713
R6138 VSS.n3437 VSS.n57 0.0147651
R6139 VSS.n3438 VSS.n54 0.0147651
R6140 VSS.n967 VSS.n966 0.0147581
R6141 VSS.n1758 VSS.n1757 0.0142813
R6142 VSS.n3340 VSS.n75 0.0140692
R6143 VSS.n3339 VSS.n3163 0.0135154
R6144 VSS.n3277 VSS.n3159 0.0135154
R6145 VSS.n1614 VSS.n1101 0.0132331
R6146 VSS.n3430 VSS.n69 0.0124077
R6147 VSS.n3358 VSS.n74 0.0124077
R6148 VSS.t191 VSS.n60 0.0121715
R6149 VSS.t319 VSS.n51 0.0121715
R6150 VSS.n3326 VSS.n3162 0.0118538
R6151 VSS.n1145 VSS.n1144 0.0115959
R6152 VSS.n3281 VSS.n3159 0.0113
R6153 VSS.n3478 VSS.n1 0.0111996
R6154 VSS.n3436 VSS.n61 0.011134
R6155 VSS.n3439 VSS.n50 0.011134
R6156 VSS.n2152 VSS.n2151 0.0110691
R6157 VSS.n2151 VSS.n613 0.0110691
R6158 VSS.n3448 VSS.n3445 0.0109186
R6159 VSS.n3428 VSS.n3427 0.0107462
R6160 VSS.n3374 VSS.n73 0.0107462
R6161 VSS.n1134 VSS.n1133 0.0106712
R6162 VSS.n3306 VSS.n3161 0.0101923
R6163 VSS.n1141 VSS.n1140 0.0100548
R6164 VSS.n1434 VSS.n1433 0.0100548
R6165 VSS.n3276 VSS.n3274 0.00978125
R6166 VSS.n3273 VSS.n3236 0.00978125
R6167 VSS.n3276 VSS.n3275 0.00969179
R6168 VSS.n3225 VSS.n3160 0.00963846
R6169 VSS.n1751 VSS.n1050 0.00959535
R6170 VSS.n1707 VSS.n1045 0.00959535
R6171 VSS.n1721 VSS.n622 0.00959535
R6172 VSS.n3173 VSS.n3165 0.00908462
R6173 VSS.n3386 VSS.n3165 0.00908462
R6174 VSS.t188 VSS.n55 0.00854035
R6175 VSS.t188 VSS.n56 0.00854035
R6176 VSS.n3293 VSS.n3160 0.00853077
R6177 VSS.n3465 VSS.n3464 0.00833133
R6178 VSS.n3466 VSS.n3465 0.00833133
R6179 VSS.n3316 VSS.n3161 0.00797692
R6180 VSS.n3447 VSS.n3446 0.00797126
R6181 VSS.n3446 VSS.t332 0.00797126
R6182 VSS.n1246 VSS.n1243 0.00782743
R6183 VSS.n1003 VSS.n1002 0.00750352
R6184 VSS.n3428 VSS.n3166 0.00742308
R6185 VSS.n3370 VSS.n73 0.00742308
R6186 VSS.n3436 VSS.t189 0.00655042
R6187 VSS.t191 VSS.n3436 0.00655042
R6188 VSS.n3437 VSS.t191 0.00655042
R6189 VSS.t188 VSS.n3437 0.00655042
R6190 VSS.n3438 VSS.t188 0.00655042
R6191 VSS.t319 VSS.n3438 0.00655042
R6192 VSS.n3439 VSS.t319 0.00655042
R6193 VSS.t190 VSS.n3439 0.00655042
R6194 VSS.n1753 VSS.n639 0.00651467
R6195 VSS.n1754 VSS.n628 0.00651467
R6196 VSS.n3207 VSS.n3162 0.00631538
R6197 VSS.n3436 VSS.n62 0.00594669
R6198 VSS.n3439 VSS.n49 0.00594669
R6199 VSS.n3431 VSS.n3430 0.00576154
R6200 VSS.n3199 VSS.n74 0.00576154
R6201 VSS.n1050 VSS.n1046 0.00554309
R6202 VSS.n1707 VSS.n1706 0.00554309
R6203 VSS.n1043 VSS.n1013 0.00554309
R6204 VSS.n1040 VSS.n1013 0.00554309
R6205 VSS.n1041 VSS.n1014 0.00554309
R6206 VSS.n1037 VSS.n1014 0.00554309
R6207 VSS.n1038 VSS.n1015 0.00554309
R6208 VSS.n1034 VSS.n1015 0.00554309
R6209 VSS.n1035 VSS.n1016 0.00554309
R6210 VSS.n1031 VSS.n1016 0.00554309
R6211 VSS.n1032 VSS.n1017 0.00554309
R6212 VSS.n1028 VSS.n1017 0.00554309
R6213 VSS.n1029 VSS.n1018 0.00554309
R6214 VSS.n1025 VSS.n1018 0.00554309
R6215 VSS.n1026 VSS.n1019 0.00554309
R6216 VSS.n1022 VSS.n1019 0.00554309
R6217 VSS.n1023 VSS.n1021 0.00554309
R6218 VSS.n1021 VSS.n1020 0.00554309
R6219 VSS.n1024 VSS.n1022 0.00554309
R6220 VSS.n1024 VSS.n1023 0.00554309
R6221 VSS.n1027 VSS.n1025 0.00554309
R6222 VSS.n1027 VSS.n1026 0.00554309
R6223 VSS.n1030 VSS.n1028 0.00554309
R6224 VSS.n1030 VSS.n1029 0.00554309
R6225 VSS.n1033 VSS.n1031 0.00554309
R6226 VSS.n1033 VSS.n1032 0.00554309
R6227 VSS.n1036 VSS.n1034 0.00554309
R6228 VSS.n1036 VSS.n1035 0.00554309
R6229 VSS.n1039 VSS.n1037 0.00554309
R6230 VSS.n1039 VSS.n1038 0.00554309
R6231 VSS.n1042 VSS.n1040 0.00554309
R6232 VSS.n1042 VSS.n1041 0.00554309
R6233 VSS.n1706 VSS.n1044 0.00554309
R6234 VSS.n1044 VSS.n1043 0.00554309
R6235 VSS.n1046 VSS.n1045 0.00554309
R6236 VSS.n1020 VSS.n627 0.00554309
R6237 VSS.n1702 VSS.n1051 0.00554309
R6238 VSS.n1748 VSS.n1736 0.00554309
R6239 VSS.n1737 VSS.n1708 0.00554309
R6240 VSS.n1735 VSS.n1734 0.00554309
R6241 VSS.n1739 VSS.n1709 0.00554309
R6242 VSS.n1733 VSS.n1732 0.00554309
R6243 VSS.n1740 VSS.n1710 0.00554309
R6244 VSS.n1731 VSS.n1730 0.00554309
R6245 VSS.n1741 VSS.n1711 0.00554309
R6246 VSS.n1729 VSS.n1728 0.00554309
R6247 VSS.n1742 VSS.n1712 0.00554309
R6248 VSS.n1727 VSS.n1726 0.00554309
R6249 VSS.n1743 VSS.n1713 0.00554309
R6250 VSS.n1725 VSS.n1724 0.00554309
R6251 VSS.n1744 VSS.n1714 0.00554309
R6252 VSS.n1723 VSS.n1722 0.00554309
R6253 VSS.n1745 VSS.n1717 0.00554309
R6254 VSS.n1721 VSS.n1718 0.00554309
R6255 VSS.n1756 VSS.n624 0.00554309
R6256 VSS.n624 VSS.n622 0.00554309
R6257 VSS.n1718 VSS.n1717 0.00554309
R6258 VSS.n1745 VSS.n1723 0.00554309
R6259 VSS.n1722 VSS.n1714 0.00554309
R6260 VSS.n1744 VSS.n1725 0.00554309
R6261 VSS.n1724 VSS.n1713 0.00554309
R6262 VSS.n1743 VSS.n1727 0.00554309
R6263 VSS.n1726 VSS.n1712 0.00554309
R6264 VSS.n1742 VSS.n1729 0.00554309
R6265 VSS.n1728 VSS.n1711 0.00554309
R6266 VSS.n1741 VSS.n1731 0.00554309
R6267 VSS.n1730 VSS.n1710 0.00554309
R6268 VSS.n1740 VSS.n1733 0.00554309
R6269 VSS.n1732 VSS.n1709 0.00554309
R6270 VSS.n1739 VSS.n1735 0.00554309
R6271 VSS.n1734 VSS.n1708 0.00554309
R6272 VSS.n1748 VSS.n1737 0.00554309
R6273 VSS.n1736 VSS.n1702 0.00554309
R6274 VSS.n1750 VSS.n1051 0.00554309
R6275 VSS.n1600 VSS.n1599 0.00508015
R6276 VSS.n1747 VSS.n1746 0.00507377
R6277 VSS.n1749 VSS.n1701 0.00507377
R6278 VSS.t191 VSS.n59 0.00490922
R6279 VSS.t319 VSS.n52 0.00490922
R6280 VSS.n3349 VSS.n3163 0.00465385
R6281 VSS.n3336 VSS.n75 0.0041
R6282 VSS.n1387 VSS.n1386 0.0041
R6283 VSS.n2210 VSS.n594 0.00405263
R6284 VSS.n617 VSS.n595 0.00405263
R6285 VSS.n1113 VSS.n1112 0.00372171
R6286 VSS.n639 VSS.n627 0.00358068
R6287 VSS.n1756 VSS.n628 0.00358068
R6288 VSS.n3445 VSS.n39 0.00338889
R6289 VSS.n39 VSS.n37 0.00338889
R6290 VSS.n1720 VSS.n1053 0.00328572
R6291 VSS.n1716 VSS.n1053 0.00328572
R6292 VSS.n1719 VSS.n1052 0.00328572
R6293 VSS.n1715 VSS.n1052 0.00328572
R6294 VSS.n1746 VSS.n1738 0.00328572
R6295 VSS.n1747 VSS.n1700 0.00328572
R6296 VSS.n1720 VSS.n1697 0.00328572
R6297 VSS.n1719 VSS.n1698 0.00328572
R6298 VSS.n1738 VSS.n1699 0.00328572
R6299 VSS.n1716 VSS.n1698 0.00328572
R6300 VSS.n1715 VSS.n1699 0.00328572
R6301 VSS.n1701 VSS.n1700 0.00328572
R6302 VSS.n1426 VSS.n1425 0.00327397
R6303 VSS.n3417 VSS.n71 0.00299231
R6304 VSS.n3189 VSS.n3164 0.00299231
R6305 VSS.n1584 VSS.n1571 0.00296575
R6306 VSS.n1047 VSS.n1008 0.00296393
R6307 VSS.n1705 VSS.n1006 0.00296393
R6308 VSS.n1048 VSS.n1009 0.00296393
R6309 VSS.n1704 VSS.n1005 0.00296393
R6310 VSS.n1049 VSS.n1010 0.00296393
R6311 VSS.n1703 VSS.n1004 0.00296393
R6312 VSS.n1752 VSS.n1011 0.00296393
R6313 VSS.n1012 VSS.n1003 0.00296393
R6314 VSS.n1705 VSS.n1008 0.00296393
R6315 VSS.n1704 VSS.n1009 0.00296393
R6316 VSS.n1703 VSS.n1010 0.00296393
R6317 VSS.n1752 VSS.n1012 0.00296393
R6318 VSS.n1047 VSS.n1007 0.00296393
R6319 VSS.n1048 VSS.n1006 0.00296393
R6320 VSS.n1049 VSS.n1005 0.00296393
R6321 VSS.n1011 VSS.n1004 0.00296393
R6322 VSS.n2153 VSS.n2152 0.00272514
R6323 VSS.n3218 VSS.n76 0.00243846
R6324 VSS.n3437 VSS.n58 0.00231556
R6325 VSS.n3438 VSS.n53 0.00231556
R6326 VSS.n2152 VSS.n1759 0.00220437
R6327 VSS.n3232 VSS.n78 0.00188462
R6328 VSS.n3396 VSS.n72 0.00133077
R6329 VSS.t189 VSS.n63 0.0012781
R6330 VSS.t190 VSS.n48 0.0012781
R6331 VSS.n1002 VSS.t338 0.00100704
R6332 VSS.n3303 VSS.n77 0.000776923
R6333 VSS.n1364 VSS.n1216 0.000659292
R6334 VDD.t262 VDD.t38 864.865
R6335 VDD.t142 VDD.n14 706.564
R6336 VDD.n14 VDD.t262 648.649
R6337 VDD.t284 VDD.t145 629.345
R6338 VDD.n394 VDD.t242 589.355
R6339 VDD.n393 VDD.t167 589.355
R6340 VDD.n400 VDD.t165 589.355
R6341 VDD.n407 VDD.t200 589.355
R6342 VDD.n414 VDD.t204 589.355
R6343 VDD.n421 VDD.t206 589.355
R6344 VDD.n428 VDD.t169 589.355
R6345 VDD.n435 VDD.t202 589.355
R6346 VDD.n30 VDD.t359 552.125
R6347 VDD.t145 VDD.t21 501.932
R6348 VDD.t154 VDD.n247 484.969
R6349 VDD.n254 VDD.t150 480.769
R6350 VDD.t363 VDD.t142 471.043
R6351 VDD.t280 VDD.t270 471.043
R6352 VDD.t285 VDD.t336 471.043
R6353 VDD.t359 VDD.t87 471.043
R6354 VDD.n261 VDD.t274 448.111
R6355 VDD.t352 VDD.n260 443.911
R6356 VDD.n260 VDD.t82 443.911
R6357 VDD.n255 VDD.t84 443.911
R6358 VDD.n255 VDD.t339 443.911
R6359 VDD.t339 VDD.n254 443.911
R6360 VDD.t21 VDD.t19 432.433
R6361 VDD.n401 VDD.t131 419.211
R6362 VDD.n408 VDD.t81 419.211
R6363 VDD.n415 VDD.t80 419.211
R6364 VDD.n422 VDD.t69 419.211
R6365 VDD.n429 VDD.t147 419.211
R6366 VDD.n436 VDD.t162 419.211
R6367 VDD.t57 VDD.t103 416.988
R6368 VDD.t208 VDD.t0 403.476
R6369 VDD.t270 VDD.t363 393.822
R6370 VDD.t336 VDD.t280 393.822
R6371 VDD.t87 VDD.t285 393.822
R6372 VDD.t313 VDD.t316 384.764
R6373 VDD.t17 VDD.t297 372.587
R6374 VDD.t311 VDD.t15 372.228
R6375 VDD.t34 VDD.t25 372.228
R6376 VDD.n30 VDD.t284 355.212
R6377 VDD.t150 VDD.t152 346.154
R6378 VDD.t152 VDD.t177 346.154
R6379 VDD.t177 VDD.t154 346.154
R6380 VDD.n514 VDD.t92 345.56
R6381 VDD.t92 VDD.t115 335.908
R6382 VDD.n515 VDD.t318 320.464
R6383 VDD.t86 VDD.t8 288.611
R6384 VDD.t13 VDD.t129 282.546
R6385 VDD.n564 VDD.t171 282.116
R6386 VDD.n528 VDD.t299 282.116
R6387 VDD.n466 VDD.t123 281.861
R6388 VDD.t54 VDD.n471 279.923
R6389 VDD.n470 VDD.t76 278.959
R6390 VDD.t215 VDD.t240 277.027
R6391 VDD.t56 VDD.t86 275.098
R6392 VDD.t274 VDD.t276 272.437
R6393 VDD.t276 VDD.t293 272.437
R6394 VDD.t293 VDD.t101 272.437
R6395 VDD.t101 VDD.t354 272.437
R6396 VDD.t354 VDD.t348 272.437
R6397 VDD.t348 VDD.t355 272.437
R6398 VDD.t355 VDD.t349 272.437
R6399 VDD.t349 VDD.t128 272.437
R6400 VDD.t128 VDD.t127 272.437
R6401 VDD.t127 VDD.t125 272.437
R6402 VDD.t125 VDD.t126 272.437
R6403 VDD.t126 VDD.t64 272.437
R6404 VDD.t64 VDD.t295 272.437
R6405 VDD.t295 VDD.t350 272.437
R6406 VDD.t350 VDD.t352 272.437
R6407 VDD.t100 VDD.t82 272.437
R6408 VDD.t315 VDD.t100 272.437
R6409 VDD.t84 VDD.t315 272.437
R6410 VDD.t115 VDD.t94 239.382
R6411 VDD.t53 VDD.t74 238.188
R6412 VDD.t221 VDD.t231 235.522
R6413 VDD.t136 VDD.t96 235.522
R6414 VDD.n542 VDD.t235 233.591
R6415 VDD.t223 VDD.t160 231.661
R6416 VDD.t51 VDD.n469 224.436
R6417 VDD.n464 VDD.t11 219.865
R6418 VDD.n475 VDD.n474 217.452
R6419 VDD.t42 VDD.t46 216.216
R6420 VDD.t309 VDD.n464 212.15
R6421 VDD.t148 VDD.t134 211.391
R6422 VDD.t8 VDD.t78 208.494
R6423 VDD.n145 VDD.n7 199.776
R6424 VDD.n147 VDD.n7 199.776
R6425 VDD.n147 VDD.n8 199.776
R6426 VDD.n145 VDD.n8 199.776
R6427 VDD.n370 VDD.n342 199.776
R6428 VDD.n370 VDD.n343 199.776
R6429 VDD.n368 VDD.n342 199.776
R6430 VDD.n368 VDD.n343 199.776
R6431 VDD.n382 VDD.n376 199.776
R6432 VDD.n382 VDD.n377 199.776
R6433 VDD.n380 VDD.n376 199.776
R6434 VDD.n380 VDD.n377 199.776
R6435 VDD.t72 VDD.t219 196.911
R6436 VDD.t23 VDD.t217 196.911
R6437 VDD.t217 VDD.t307 196.911
R6438 VDD.t181 VDD.t305 196.911
R6439 VDD.t328 VDD.t60 196.911
R6440 VDD.t103 VDD.t208 196.911
R6441 VDD.t225 VDD.t229 196.911
R6442 VDD.t330 VDD.t65 196.721
R6443 VDD.t334 VDD.t70 196.721
R6444 VDD.t27 VDD.t109 196.721
R6445 VDD.t279 VDD.n145 187.815
R6446 VDD.n147 VDD.t141 187.815
R6447 VDD.n370 VDD.t111 187.815
R6448 VDD.t238 VDD.n368 187.815
R6449 VDD.n382 VDD.t320 187.815
R6450 VDD.t266 VDD.n380 187.815
R6451 VDD.t289 VDD.t44 181.468
R6452 VDD.t175 VDD.t328 174.71
R6453 VDD.t109 VDD.t260 174.542
R6454 VDD.t29 VDD.t227 173.745
R6455 VDD.t305 VDD.t175 168.919
R6456 VDD.t260 VDD.t334 168.756
R6457 VDD.t303 VDD.t2 167.954
R6458 VDD.t96 VDD.t120 167.954
R6459 VDD.t49 VDD.t42 166.024
R6460 VDD.t332 VDD.t98 162.162
R6461 VDD.n443 VDD.t36 156.802
R6462 VDD.t291 VDD.t215 155.405
R6463 VDD.n471 VDD.t303 152.511
R6464 VDD.t94 VDD.t56 150.579
R6465 VDD.t4 VDD.t48 150.579
R6466 VDD.t301 VDD.t330 149.47
R6467 VDD.t356 VDD.t13 149.47
R6468 VDD.t78 VDD.t102 142.857
R6469 VDD.t32 VDD.t278 142.857
R6470 VDD.n513 VDD.t57 138.031
R6471 VDD.t229 VDD.t287 121.623
R6472 VDD.t235 VDD.t6 119.692
R6473 VDD.t67 VDD.t158 119.692
R6474 VDD.t287 VDD.t233 113.9
R6475 VDD.t2 VDD.n470 111.969
R6476 VDD.t122 VDD.t279 107.053
R6477 VDD.t282 VDD.t122 107.053
R6478 VDD.t114 VDD.t282 107.053
R6479 VDD.t268 VDD.t114 107.053
R6480 VDD.t327 VDD.t268 107.053
R6481 VDD.t89 VDD.t327 107.053
R6482 VDD.t63 VDD.t89 107.053
R6483 VDD.t366 VDD.t63 107.053
R6484 VDD.t338 VDD.t366 107.053
R6485 VDD.t113 VDD.t144 107.053
R6486 VDD.t362 VDD.t113 107.053
R6487 VDD.t361 VDD.t362 107.053
R6488 VDD.t62 VDD.t361 107.053
R6489 VDD.t365 VDD.t62 107.053
R6490 VDD.t283 VDD.t365 107.053
R6491 VDD.t269 VDD.t283 107.053
R6492 VDD.t112 VDD.t269 107.053
R6493 VDD.t141 VDD.t112 107.053
R6494 VDD.t111 VDD.t343 107.053
R6495 VDD.t343 VDD.t272 107.053
R6496 VDD.t272 VDD.t264 107.053
R6497 VDD.t264 VDD.t118 107.053
R6498 VDD.t118 VDD.t117 107.053
R6499 VDD.t117 VDD.t105 107.053
R6500 VDD.t105 VDD.t325 107.053
R6501 VDD.t325 VDD.t324 107.053
R6502 VDD.t324 VDD.t273 107.053
R6503 VDD.t183 VDD.t265 107.053
R6504 VDD.t265 VDD.t239 107.053
R6505 VDD.t239 VDD.t197 107.053
R6506 VDD.t197 VDD.t196 107.053
R6507 VDD.t196 VDD.t326 107.053
R6508 VDD.t326 VDD.t342 107.053
R6509 VDD.t342 VDD.t185 107.053
R6510 VDD.t185 VDD.t184 107.053
R6511 VDD.t184 VDD.t238 107.053
R6512 VDD.t320 VDD.t321 107.053
R6513 VDD.t321 VDD.t149 107.053
R6514 VDD.t149 VDD.t195 107.053
R6515 VDD.t195 VDD.t108 107.053
R6516 VDD.t108 VDD.t199 107.053
R6517 VDD.t199 VDD.t187 107.053
R6518 VDD.t187 VDD.t322 107.053
R6519 VDD.t322 VDD.t267 107.053
R6520 VDD.t267 VDD.t106 107.053
R6521 VDD.t341 VDD.t107 107.053
R6522 VDD.t107 VDD.t237 107.053
R6523 VDD.t237 VDD.t344 107.053
R6524 VDD.t344 VDD.t194 107.053
R6525 VDD.t194 VDD.t138 107.053
R6526 VDD.t138 VDD.t198 107.053
R6527 VDD.t198 VDD.t186 107.053
R6528 VDD.t186 VDD.t323 107.053
R6529 VDD.t323 VDD.t266 107.053
R6530 VDD.t36 VDD.t53 98.3612
R6531 VDD.t158 VDD.t32 88.8036
R6532 VDD.n541 VDD.t40 87.8383
R6533 VDD.t65 VDD.t311 85.825
R6534 VDD.t6 VDD.t221 77.2206
R6535 VDD.t134 VDD.t67 77.2206
R6536 VDD.t102 VDD.n513 71.4291
R6537 VDD.t132 VDD.n541 67.5681
R6538 VDD.n189 VDD.n188 66.6672
R6539 VDD.n201 VDD.n175 66.6672
R6540 VDD.n203 VDD.n202 66.6672
R6541 VDD.n215 VDD.n167 66.6672
R6542 VDD.n217 VDD.n216 66.6672
R6543 VDD.n230 VDD.n159 66.6672
R6544 VDD.n232 VDD.n231 66.6672
R6545 VDD.t240 VDD.t181 66.6028
R6546 VDD.n329 VDD.n328 66.5439
R6547 VDD.n327 VDD.n282 66.5439
R6548 VDD.n319 VDD.n318 66.5439
R6549 VDD.n317 VDD.n286 66.5439
R6550 VDD.n309 VDD.n308 66.5439
R6551 VDD.n307 VDD.n290 66.5439
R6552 VDD.n299 VDD.n298 66.5439
R6553 VDD.t70 VDD.t309 66.5386
R6554 VDD.t252 VDD.n187 66.177
R6555 VDD.t188 VDD.n279 66.0664
R6556 VDD.t227 VDD.t4 65.6376
R6557 VDD.n353 VDD.n351 65.4873
R6558 VDD.n356 VDD.n350 65.4873
R6559 VDD.t60 VDD.t17 60.8113
R6560 VDD.t129 VDD.t27 60.7527
R6561 VDD.n189 VDD.t173 59.877
R6562 VDD.t256 VDD.n201 59.877
R6563 VDD.n203 VDD.t213 59.877
R6564 VDD.t244 VDD.n215 59.877
R6565 VDD.n217 VDD.t156 59.877
R6566 VDD.t211 VDD.n230 59.877
R6567 VDD.n232 VDD.t254 59.877
R6568 VDD.t297 VDD.t51 59.8461
R6569 VDD.t15 VDD.t34 59.7883
R6570 VDD.t25 VDD.t11 59.7883
R6571 VDD.n328 VDD.t248 59.7664
R6572 VDD.t192 VDD.n282 59.7664
R6573 VDD.n318 VDD.t258 59.7664
R6574 VDD.t190 VDD.n286 59.7664
R6575 VDD.n308 VDD.t179 59.7664
R6576 VDD.t246 VDD.n290 59.7664
R6577 VDD.n298 VDD.t250 59.7664
R6578 VDD.n474 VDD.t72 56.9503
R6579 VDD.n146 VDD.t338 53.527
R6580 VDD.t144 VDD.n146 53.527
R6581 VDD.t273 VDD.n369 53.527
R6582 VDD.n369 VDD.t183 53.527
R6583 VDD.t106 VDD.n381 53.527
R6584 VDD.n381 VDD.t341 53.527
R6585 VDD.t40 VDD.t49 50.1936
R6586 VDD.t0 VDD.t299 48.263
R6587 VDD.t120 VDD.t171 48.263
R6588 VDD.t123 VDD.t313 48.2165
R6589 VDD.n354 VDD.n350 48.0418
R6590 VDD.n355 VDD.n351 48.0418
R6591 VDD.t74 VDD.t301 47.2522
R6592 VDD.t316 VDD.t356 47.2522
R6593 VDD.n475 VDD.t163 44.4358
R6594 VDD.t76 VDD.t291 41.5063
R6595 VDD.t219 VDD.t332 34.7495
R6596 VDD.t98 VDD.t23 34.7495
R6597 VDD.t46 VDD.t289 34.7495
R6598 VDD.t307 VDD.t54 29.9233
R6599 VDD.t160 VDD.t148 24.1318
R6600 VDD.t231 VDD.t29 23.1665
R6601 VDD.n522 VDD.t90 21.6375
R6602 VDD.n522 VDD.t58 21.6375
R6603 VDD.n556 VDD.t50 21.6375
R6604 VDD.t48 VDD.t223 19.3055
R6605 VDD.n541 VDD.t10 16.2012
R6606 VDD.n513 VDD.t59 15.981
R6607 VDD.t44 VDD.t136 15.4445
R6608 VDD.n246 VDD.t340 12.2195
R6609 VDD.n235 VDD.t254 12.1776
R6610 VDD.t250 VDD.n297 12.1637
R6611 VDD.n236 VDD.n235 11.4951
R6612 VDD.n297 VDD.n294 11.4938
R6613 VDD.n254 VDD.n253 11.0111
R6614 VDD.n256 VDD.n255 11.0111
R6615 VDD.n260 VDD.n259 11.0111
R6616 VDD.n257 VDD.t85 10.0145
R6617 VDD.n258 VDD.t83 10.0145
R6618 VDD.n245 VDD.t353 10.0145
R6619 VDD.n567 VDD.n150 9.48313
R6620 VDD.n249 VDD.t155 9.42355
R6621 VDD.n252 VDD.t151 9.42355
R6622 VDD.n244 VDD.n243 8.54446
R6623 VDD.n242 VDD.n241 8.54446
R6624 VDD.n394 VDD.t243 8.52192
R6625 VDD.n393 VDD.t168 8.52192
R6626 VDD.n400 VDD.t166 8.46717
R6627 VDD.n407 VDD.t201 8.46717
R6628 VDD.n414 VDD.t205 8.46717
R6629 VDD.n421 VDD.t207 8.46717
R6630 VDD.n428 VDD.t170 8.46717
R6631 VDD.n435 VDD.t203 8.46717
R6632 VDD.n251 VDD.n250 8.11105
R6633 VDD.n515 VDD.n514 7.72251
R6634 VDD.n562 VDD.t172 7.51784
R6635 VDD.n554 VDD.t133 7.5061
R6636 VDD.n479 VDD.t333 7.46
R6637 VDD.n482 VDD.t308 7.46
R6638 VDD.n512 VDD.t95 7.40883
R6639 VDD.n511 VDD.t346 7.40883
R6640 VDD.n538 VDD.t5 7.40883
R6641 VDD.n35 VDD.t20 6.91104
R6642 VDD.n188 VDD.t252 6.79062
R6643 VDD.t173 VDD.n175 6.79062
R6644 VDD.n202 VDD.t256 6.79062
R6645 VDD.t213 VDD.n167 6.79062
R6646 VDD.n216 VDD.t244 6.79062
R6647 VDD.t156 VDD.n159 6.79062
R6648 VDD.n231 VDD.t211 6.79062
R6649 VDD.n329 VDD.t188 6.77807
R6650 VDD.t248 VDD.n327 6.77807
R6651 VDD.n319 VDD.t192 6.77807
R6652 VDD.t258 VDD.n317 6.77807
R6653 VDD.n309 VDD.t190 6.77807
R6654 VDD.t179 VDD.n307 6.77807
R6655 VDD.n299 VDD.t246 6.77807
R6656 VDD.n234 VDD.n155 6.3005
R6657 VDD.n233 VDD.n158 6.3005
R6658 VDD.n233 VDD.n232 6.3005
R6659 VDD.n163 VDD.n156 6.3005
R6660 VDD.n231 VDD.n156 6.3005
R6661 VDD.n229 VDD.n228 6.3005
R6662 VDD.n230 VDD.n229 6.3005
R6663 VDD.n221 VDD.n160 6.3005
R6664 VDD.n160 VDD.n159 6.3005
R6665 VDD.n219 VDD.n218 6.3005
R6666 VDD.n218 VDD.n217 6.3005
R6667 VDD.n171 VDD.n166 6.3005
R6668 VDD.n216 VDD.n166 6.3005
R6669 VDD.n214 VDD.n213 6.3005
R6670 VDD.n215 VDD.n214 6.3005
R6671 VDD.n207 VDD.n168 6.3005
R6672 VDD.n168 VDD.n167 6.3005
R6673 VDD.n205 VDD.n204 6.3005
R6674 VDD.n204 VDD.n203 6.3005
R6675 VDD.n179 VDD.n174 6.3005
R6676 VDD.n202 VDD.n174 6.3005
R6677 VDD.n200 VDD.n199 6.3005
R6678 VDD.n201 VDD.n200 6.3005
R6679 VDD.n193 VDD.n176 6.3005
R6680 VDD.n176 VDD.n175 6.3005
R6681 VDD.n191 VDD.n190 6.3005
R6682 VDD.n190 VDD.n189 6.3005
R6683 VDD.n183 VDD.n182 6.3005
R6684 VDD.n188 VDD.n182 6.3005
R6685 VDD.n187 VDD.n186 6.3005
R6686 VDD.n279 VDD.n278 6.3005
R6687 VDD.n331 VDD.n330 6.3005
R6688 VDD.n330 VDD.n329 6.3005
R6689 VDD.n281 VDD.n280 6.3005
R6690 VDD.n328 VDD.n281 6.3005
R6691 VDD.n326 VDD.n325 6.3005
R6692 VDD.n327 VDD.n326 6.3005
R6693 VDD.n324 VDD.n323 6.3005
R6694 VDD.n324 VDD.n282 6.3005
R6695 VDD.n320 VDD.n285 6.3005
R6696 VDD.n320 VDD.n319 6.3005
R6697 VDD.n284 VDD.n283 6.3005
R6698 VDD.n318 VDD.n284 6.3005
R6699 VDD.n316 VDD.n315 6.3005
R6700 VDD.n317 VDD.n316 6.3005
R6701 VDD.n314 VDD.n313 6.3005
R6702 VDD.n314 VDD.n286 6.3005
R6703 VDD.n310 VDD.n289 6.3005
R6704 VDD.n310 VDD.n309 6.3005
R6705 VDD.n288 VDD.n287 6.3005
R6706 VDD.n308 VDD.n288 6.3005
R6707 VDD.n306 VDD.n305 6.3005
R6708 VDD.n307 VDD.n306 6.3005
R6709 VDD.n304 VDD.n303 6.3005
R6710 VDD.n304 VDD.n290 6.3005
R6711 VDD.n300 VDD.n293 6.3005
R6712 VDD.n300 VDD.n299 6.3005
R6713 VDD.n292 VDD.n291 6.3005
R6714 VDD.n298 VDD.n292 6.3005
R6715 VDD.n296 VDD.n295 6.3005
R6716 VDD.n510 VDD.t79 6.22272
R6717 VDD.n509 VDD.t91 6.22272
R6718 VDD.n535 VDD.t33 6.22272
R6719 VDD.n396 VDD.n150 6.1835
R6720 VDD.n392 VDD.n150 6.09991
R6721 VDD.n187 VDD.n182 6.0755
R6722 VDD.n190 VDD.n182 6.0755
R6723 VDD.n190 VDD.n176 6.0755
R6724 VDD.n200 VDD.n176 6.0755
R6725 VDD.n200 VDD.n174 6.0755
R6726 VDD.n204 VDD.n174 6.0755
R6727 VDD.n204 VDD.n168 6.0755
R6728 VDD.n214 VDD.n168 6.0755
R6729 VDD.n214 VDD.n166 6.0755
R6730 VDD.n218 VDD.n166 6.0755
R6731 VDD.n218 VDD.n160 6.0755
R6732 VDD.n229 VDD.n160 6.0755
R6733 VDD.n229 VDD.n156 6.0755
R6734 VDD.n233 VDD.n156 6.0755
R6735 VDD.n234 VDD.n233 6.0755
R6736 VDD.n330 VDD.n279 6.0755
R6737 VDD.n330 VDD.n281 6.0755
R6738 VDD.n326 VDD.n281 6.0755
R6739 VDD.n326 VDD.n324 6.0755
R6740 VDD.n324 VDD.n320 6.0755
R6741 VDD.n320 VDD.n284 6.0755
R6742 VDD.n316 VDD.n284 6.0755
R6743 VDD.n316 VDD.n314 6.0755
R6744 VDD.n314 VDD.n310 6.0755
R6745 VDD.n310 VDD.n288 6.0755
R6746 VDD.n306 VDD.n288 6.0755
R6747 VDD.n306 VDD.n304 6.0755
R6748 VDD.n304 VDD.n300 6.0755
R6749 VDD.n300 VDD.n292 6.0755
R6750 VDD.n296 VDD.n292 6.0755
R6751 VDD.n520 VDD.n511 5.49789
R6752 VDD.n520 VDD.n512 5.49789
R6753 VDD.n550 VDD.n538 5.49789
R6754 VDD.n521 VDD.n509 5.41359
R6755 VDD.n521 VDD.n510 5.41359
R6756 VDD.n553 VDD.n535 5.41359
R6757 VDD.n56 VDD.n25 5.39615
R6758 VDD.n64 VDD.n22 5.39615
R6759 VDD.n71 VDD.n19 5.39615
R6760 VDD.n557 VDD.n534 5.35702
R6761 VDD.n552 VDD.n536 5.35702
R6762 VDD.n549 VDD.n539 5.35702
R6763 VDD.n547 VDD.n540 5.35702
R6764 VDD.n545 VDD.n543 5.35702
R6765 VDD.n523 VDD.n507 5.35271
R6766 VDD.n523 VDD.n508 5.35271
R6767 VDD.n558 VDD.n533 5.35271
R6768 VDD.n559 VDD.n532 5.31398
R6769 VDD.n36 VDD.n34 5.30638
R6770 VDD.n481 VDD.n472 5.30615
R6771 VDD.n478 VDD.n473 5.29976
R6772 VDD.n445 VDD.n442 5.29976
R6773 VDD.n551 VDD.n537 5.28659
R6774 VDD.n510 VDD.t9 5.05606
R6775 VDD.n509 VDD.t31 5.05606
R6776 VDD.n535 VDD.t68 5.05606
R6777 VDD.n374 VDD.n373 4.94375
R6778 VDD.n480 VDD.t99 4.70061
R6779 VDD.n447 VDD.t66 4.70061
R6780 VDD.n185 VDD.n184 4.60502
R6781 VDD.n247 VDD.n153 4.56013
R6782 VDD.n247 VDD.n151 4.56013
R6783 VDD.n249 VDD.n248 4.55193
R6784 VDD.n402 VDD.n399 4.5005
R6785 VDD.n399 VDD.n398 4.5005
R6786 VDD.n402 VDD.n401 4.5005
R6787 VDD.n401 VDD.n398 4.5005
R6788 VDD.n409 VDD.n406 4.5005
R6789 VDD.n406 VDD.n405 4.5005
R6790 VDD.n409 VDD.n408 4.5005
R6791 VDD.n408 VDD.n405 4.5005
R6792 VDD.n416 VDD.n413 4.5005
R6793 VDD.n413 VDD.n412 4.5005
R6794 VDD.n416 VDD.n415 4.5005
R6795 VDD.n415 VDD.n412 4.5005
R6796 VDD.n423 VDD.n420 4.5005
R6797 VDD.n420 VDD.n419 4.5005
R6798 VDD.n423 VDD.n422 4.5005
R6799 VDD.n422 VDD.n419 4.5005
R6800 VDD.n430 VDD.n427 4.5005
R6801 VDD.n427 VDD.n426 4.5005
R6802 VDD.n430 VDD.n429 4.5005
R6803 VDD.n429 VDD.n426 4.5005
R6804 VDD.n437 VDD.n434 4.5005
R6805 VDD.n434 VDD.n433 4.5005
R6806 VDD.n437 VDD.n436 4.5005
R6807 VDD.n436 VDD.n433 4.5005
R6808 VDD.n238 VDD.n237 4.5005
R6809 VDD.n157 VDD.n154 4.5005
R6810 VDD.n225 VDD.n224 4.5005
R6811 VDD.n227 VDD.n226 4.5005
R6812 VDD.n223 VDD.n222 4.5005
R6813 VDD.n220 VDD.n164 4.5005
R6814 VDD.n210 VDD.n165 4.5005
R6815 VDD.n212 VDD.n211 4.5005
R6816 VDD.n209 VDD.n208 4.5005
R6817 VDD.n206 VDD.n172 4.5005
R6818 VDD.n196 VDD.n173 4.5005
R6819 VDD.n198 VDD.n197 4.5005
R6820 VDD.n195 VDD.n194 4.5005
R6821 VDD.n192 VDD.n180 4.5005
R6822 VDD.n184 VDD.n181 4.5005
R6823 VDD.n467 VDD.n441 4.5005
R6824 VDD.n333 VDD.n270 4.5005
R6825 VDD.n333 VDD.n271 4.5005
R6826 VDD.n333 VDD.n269 4.5005
R6827 VDD.n333 VDD.n272 4.5005
R6828 VDD.n333 VDD.n268 4.5005
R6829 VDD.n333 VDD.n273 4.5005
R6830 VDD.n333 VDD.n267 4.5005
R6831 VDD.n333 VDD.n274 4.5005
R6832 VDD.n333 VDD.n266 4.5005
R6833 VDD.n333 VDD.n275 4.5005
R6834 VDD.n333 VDD.n265 4.5005
R6835 VDD.n333 VDD.n276 4.5005
R6836 VDD.n333 VDD.n264 4.5005
R6837 VDD.n333 VDD.n277 4.5005
R6838 VDD.n333 VDD.n263 4.5005
R6839 VDD.n333 VDD.n332 4.5005
R6840 VDD.n360 VDD.n359 4.5005
R6841 VDD.n366 VDD.n365 4.5005
R6842 VDD.n364 VDD.n346 4.5005
R6843 VDD.n363 VDD.n362 4.5005
R6844 VDD.n361 VDD.n347 4.5005
R6845 VDD.n389 VDD.n337 4.5005
R6846 VDD.n388 VDD.n387 4.5005
R6847 VDD.n386 VDD.n339 4.5005
R6848 VDD.n385 VDD.n384 4.5005
R6849 VDD.n391 VDD.n390 4.5005
R6850 VDD.n496 VDD.t61 4.46351
R6851 VDD.n494 VDD.t329 4.46351
R6852 VDD.n493 VDD.t306 4.46351
R6853 VDD.n491 VDD.t182 4.46351
R6854 VDD.n490 VDD.t216 4.46351
R6855 VDD.n488 VDD.t77 4.46351
R6856 VDD.n453 VDD.t317 4.46351
R6857 VDD.n455 VDD.t14 4.46351
R6858 VDD.n456 VDD.t28 4.46351
R6859 VDD.n458 VDD.t110 4.46351
R6860 VDD.n459 VDD.t335 4.46351
R6861 VDD.n461 VDD.t71 4.46351
R6862 VDD.n516 VDD.t345 4.45405
R6863 VDD.n544 VDD.t234 4.385
R6864 VDD.n499 VDD.t298 4.36426
R6865 VDD.n485 VDD.t304 4.36426
R6866 VDD.n483 VDD.t55 4.36426
R6867 VDD.n476 VDD.t164 4.36426
R6868 VDD.n526 VDD.t300 4.36426
R6869 VDD.n465 VDD.t124 4.36426
R6870 VDD.n451 VDD.t26 4.36426
R6871 VDD.n449 VDD.t16 4.36426
R6872 VDD.n443 VDD.t37 4.36426
R6873 VDD.n487 VDD.t3 4.36035
R6874 VDD.n489 VDD.t292 4.36035
R6875 VDD.n492 VDD.t241 4.36035
R6876 VDD.n495 VDD.t176 4.36035
R6877 VDD.n497 VDD.t18 4.36035
R6878 VDD.n501 VDD.t52 4.36035
R6879 VDD.n516 VDD.t319 4.36035
R6880 VDD.n524 VDD.t1 4.36035
R6881 VDD.n544 VDD.t288 4.36035
R6882 VDD.n560 VDD.t121 4.36035
R6883 VDD.n444 VDD.t302 4.36035
R6884 VDD.n446 VDD.t312 4.36035
R6885 VDD.n448 VDD.t35 4.36035
R6886 VDD.n450 VDD.t12 4.36035
R6887 VDD.n462 VDD.t310 4.36035
R6888 VDD.n460 VDD.t261 4.36035
R6889 VDD.n457 VDD.t130 4.36035
R6890 VDD.n454 VDD.t357 4.36035
R6891 VDD.n452 VDD.t314 4.36035
R6892 VDD.n86 VDD.t263 4.36035
R6893 VDD.n10 VDD.t39 4.36035
R6894 VDD.n486 VDD.n470 4.35926
R6895 VDD.n518 VDD.n514 4.35926
R6896 VDD.n464 VDD.n463 4.35926
R6897 VDD.n477 VDD.n474 4.35925
R6898 VDD.n484 VDD.n471 4.35925
R6899 VDD.n517 VDD.n515 4.35925
R6900 VDD.n546 VDD.n542 4.35925
R6901 VDD.n84 VDD.n14 4.35924
R6902 VDD.n31 VDD.n30 4.35914
R6903 VDD.n49 VDD.t360 4.31143
R6904 VDD.n78 VDD.t143 4.31143
R6905 VDD.n519 VDD.t93 4.29774
R6906 VDD.n519 VDD.t347 4.29774
R6907 VDD.n548 VDD.t7 4.29774
R6908 VDD.n555 VDD.t41 4.28209
R6909 VDD.n359 VDD.n358 4.1815
R6910 VDD.n532 VDD.t45 3.91054
R6911 VDD.t278 VDD.t132 3.8615
R6912 VDD.n537 VDD.t161 3.7566
R6913 VDD.n240 VDD.t275 3.20383
R6914 VDD.n476 VDD.n475 3.05229
R6915 VDD.n467 VDD.n440 2.97032
R6916 VDD.n148 VDD.n6 2.85445
R6917 VDD.n379 VDD.n378 2.85445
R6918 VDD.n379 VDD.n338 2.85445
R6919 VDD.n144 VDD.n6 2.82271
R6920 VDD.n440 VDD.n151 2.82015
R6921 VDD.n34 VDD.t146 2.81423
R6922 VDD.n404 VDD.n403 2.70462
R6923 VDD.n411 VDD.n410 2.70462
R6924 VDD.n418 VDD.n417 2.70462
R6925 VDD.n425 VDD.n424 2.70462
R6926 VDD.n432 VDD.n431 2.70462
R6927 VDD.n439 VDD.n438 2.70462
R6928 VDD.n345 VDD.n344 2.5272
R6929 VDD.n344 VDD.n340 2.5272
R6930 VDD.n372 VDD.n341 2.5272
R6931 VDD.n378 VDD.n375 2.5272
R6932 VDD.n242 VDD.n239 2.38212
R6933 VDD.n503 VDD.n469 2.29149
R6934 VDD.n360 VDD.n341 2.28609
R6935 VDD.n390 VDD.n338 2.28609
R6936 VDD.n498 VDD.n468 2.28317
R6937 VDD.n525 VDD.n506 2.28317
R6938 VDD.n561 VDD.n531 2.28317
R6939 VDD.n34 VDD.t22 2.28216
R6940 VDD.n512 VDD.t116 2.2755
R6941 VDD.n511 VDD.t119 2.2755
R6942 VDD.n538 VDD.t30 2.2755
R6943 VDD.n396 VDD.n395 2.25109
R6944 VDD.n503 VDD.n502 2.2505
R6945 VDD.n500 VDD.n468 2.2505
R6946 VDD.n527 VDD.n506 2.2505
R6947 VDD.n563 VDD.n531 2.2505
R6948 VDD.n262 VDD.n261 2.2505
R6949 VDD.n240 VDD.n152 2.2505
R6950 VDD.n37 VDD.n33 2.2505
R6951 VDD.n39 VDD.n38 2.2505
R6952 VDD.n40 VDD.n32 2.2505
R6953 VDD.n42 VDD.n41 2.2505
R6954 VDD.n43 VDD.n29 2.2505
R6955 VDD.n45 VDD.n44 2.2505
R6956 VDD.n46 VDD.n28 2.2505
R6957 VDD.n48 VDD.n47 2.2505
R6958 VDD.n50 VDD.n27 2.2505
R6959 VDD.n52 VDD.n51 2.2505
R6960 VDD.n53 VDD.n26 2.2505
R6961 VDD.n55 VDD.n54 2.2505
R6962 VDD.n57 VDD.n24 2.2505
R6963 VDD.n59 VDD.n58 2.2505
R6964 VDD.n60 VDD.n23 2.2505
R6965 VDD.n62 VDD.n61 2.2505
R6966 VDD.n63 VDD.n21 2.2505
R6967 VDD.n66 VDD.n65 2.2505
R6968 VDD.n67 VDD.n20 2.2505
R6969 VDD.n69 VDD.n68 2.2505
R6970 VDD.n70 VDD.n18 2.2505
R6971 VDD.n73 VDD.n72 2.2505
R6972 VDD.n74 VDD.n17 2.2505
R6973 VDD.n76 VDD.n75 2.2505
R6974 VDD.n77 VDD.n16 2.2505
R6975 VDD.n80 VDD.n79 2.2505
R6976 VDD.n81 VDD.n15 2.2505
R6977 VDD.n83 VDD.n82 2.2505
R6978 VDD.n85 VDD.n13 2.2505
R6979 VDD.n88 VDD.n87 2.2505
R6980 VDD.n89 VDD.n12 2.2505
R6981 VDD.n91 VDD.n90 2.2505
R6982 VDD.n92 VDD.n11 2.2505
R6983 VDD.n94 VDD.n93 2.2505
R6984 VDD.n568 VDD.n149 2.2505
R6985 VDD.n570 VDD.n569 2.2505
R6986 VDD.n571 VDD.n5 2.2505
R6987 VDD.n573 VDD.n572 2.2505
R6988 VDD.n574 VDD.n4 2.2505
R6989 VDD.n576 VDD.n575 2.2505
R6990 VDD.n577 VDD.n3 2.2505
R6991 VDD.n579 VDD.n578 2.2505
R6992 VDD.n580 VDD.n2 2.2505
R6993 VDD.n582 VDD.n581 2.2505
R6994 VDD.n584 VDD.n583 2.2505
R6995 VDD.n1 VDD.n0 2.2505
R6996 VDD.n108 VDD.n107 2.2505
R6997 VDD.n110 VDD.n109 2.2505
R6998 VDD.n111 VDD.n106 2.2505
R6999 VDD.n113 VDD.n112 2.2505
R7000 VDD.n114 VDD.n104 2.2505
R7001 VDD.n116 VDD.n115 2.2505
R7002 VDD.n117 VDD.n103 2.2505
R7003 VDD.n119 VDD.n118 2.2505
R7004 VDD.n120 VDD.n102 2.2505
R7005 VDD.n122 VDD.n121 2.2505
R7006 VDD.n123 VDD.n101 2.2505
R7007 VDD.n125 VDD.n124 2.2505
R7008 VDD.n126 VDD.n100 2.2505
R7009 VDD.n128 VDD.n127 2.2505
R7010 VDD.n129 VDD.n99 2.2505
R7011 VDD.n131 VDD.n130 2.2505
R7012 VDD.n132 VDD.n98 2.2505
R7013 VDD.n134 VDD.n133 2.2505
R7014 VDD.n135 VDD.n97 2.2505
R7015 VDD.n137 VDD.n136 2.2505
R7016 VDD.n138 VDD.n96 2.2505
R7017 VDD.n140 VDD.n139 2.2505
R7018 VDD.n141 VDD.n9 2.2505
R7019 VDD.n143 VDD.n142 2.2505
R7020 VDD.n568 VDD.n567 2.23866
R7021 VDD.n532 VDD.t97 2.22001
R7022 VDD.n536 VDD.t135 2.22001
R7023 VDD.n536 VDD.t159 2.22001
R7024 VDD.n472 VDD.t24 2.15435
R7025 VDD.n472 VDD.t218 2.15435
R7026 VDD.n508 VDD.t104 2.10455
R7027 VDD.n508 VDD.t209 2.10455
R7028 VDD.n507 VDD.t358 2.10455
R7029 VDD.n507 VDD.t210 2.10455
R7030 VDD.n533 VDD.t290 2.10455
R7031 VDD.n533 VDD.t137 2.10455
R7032 VDD.n534 VDD.t43 2.06607
R7033 VDD.n278 VDD.t189 2.04514
R7034 VDD.n186 VDD.t253 2.04159
R7035 VDD.n392 VDD.n391 2.02679
R7036 VDD.n294 VDD.t251 2.02385
R7037 VDD.n349 VDD.t140 2.0205
R7038 VDD.n236 VDD.t255 2.0203
R7039 VDD.n542 VDD.t225 1.931
R7040 VDD.n397 VDD.n392 1.88697
R7041 VDD.n142 VDD.n95 1.86758
R7042 VDD.n473 VDD.t73 1.84822
R7043 VDD.n473 VDD.t220 1.84822
R7044 VDD.n442 VDD.t75 1.84822
R7045 VDD.n442 VDD.t331 1.84822
R7046 VDD.n397 VDD.n396 1.81813
R7047 VDD.n537 VDD.t224 1.67844
R7048 VDD.n357 VDD.n356 1.5755
R7049 VDD.n353 VDD.n352 1.5755
R7050 VDD.n534 VDD.t47 1.4923
R7051 VDD.n539 VDD.t232 1.4923
R7052 VDD.n539 VDD.t228 1.4923
R7053 VDD.n540 VDD.t236 1.4923
R7054 VDD.n540 VDD.t222 1.4923
R7055 VDD.n543 VDD.t230 1.4923
R7056 VDD.n543 VDD.t226 1.4923
R7057 VDD.n25 VDD.t286 1.4923
R7058 VDD.n25 VDD.t88 1.4923
R7059 VDD.n22 VDD.t281 1.4923
R7060 VDD.n22 VDD.t337 1.4923
R7061 VDD.n19 VDD.t364 1.4923
R7062 VDD.n19 VDD.t271 1.4923
R7063 VDD.n467 VDD.n466 1.48949
R7064 VDD.n302 VDD.n301 1.47853
R7065 VDD.n312 VDD.n311 1.47853
R7066 VDD.n322 VDD.n321 1.47853
R7067 VDD.n178 VDD.n177 1.47497
R7068 VDD.n170 VDD.n169 1.47497
R7069 VDD.n162 VDD.n161 1.47497
R7070 VDD.n505 VDD.n467 1.46788
R7071 VDD.n439 VDD.n432 1.4375
R7072 VDD.n432 VDD.n425 1.4375
R7073 VDD.n425 VDD.n418 1.4375
R7074 VDD.n418 VDD.n411 1.4375
R7075 VDD.n411 VDD.n404 1.4375
R7076 VDD.n404 VDD.n397 1.4375
R7077 VDD.n355 VDD.t139 1.15641
R7078 VDD.t139 VDD.n354 1.15641
R7079 VDD.n529 VDD.n528 1.14644
R7080 VDD.n565 VDD.n564 1.14644
R7081 VDD.n334 VDD.n262 1.0851
R7082 VDD.n365 VDD.n345 1.06648
R7083 VDD.n373 VDD.n340 1.00685
R7084 VDD.n373 VDD.n372 1.00685
R7085 VDD.n375 VDD.n374 1.00685
R7086 VDD.n352 VDD.n348 0.936026
R7087 VDD.n567 VDD.n566 0.92
R7088 VDD.n243 VDD.t296 0.9105
R7089 VDD.n243 VDD.t351 0.9105
R7090 VDD.n241 VDD.t277 0.9105
R7091 VDD.n241 VDD.t294 0.9105
R7092 VDD.n250 VDD.t153 0.813
R7093 VDD.n250 VDD.t178 0.813
R7094 VDD.n95 VDD.n10 0.791847
R7095 VDD.n145 VDD.n144 0.788
R7096 VDD.n148 VDD.n147 0.788
R7097 VDD.n350 VDD.n349 0.788
R7098 VDD.n351 VDD.n348 0.788
R7099 VDD.n368 VDD.n367 0.788
R7100 VDD.n371 VDD.n370 0.788
R7101 VDD.n380 VDD.n379 0.788
R7102 VDD.n383 VDD.n382 0.788
R7103 VDD.n335 VDD.n238 0.7505
R7104 VDD.n357 VDD.n349 0.734526
R7105 VDD.n352 VDD.n349 0.734526
R7106 VDD.n358 VDD.n348 0.676711
R7107 VDD.n244 VDD.n242 0.656214
R7108 VDD.n149 VDD.n148 0.607041
R7109 VDD.n144 VDD.n143 0.576984
R7110 VDD.n566 VDD.n565 0.563
R7111 VDD.n530 VDD.n529 0.563
R7112 VDD.n505 VDD.n504 0.563
R7113 VDD.n336 VDD.n152 0.557449
R7114 VDD.n335 VDD.n334 0.54104
R7115 VDD.n35 VDD.n33 0.511015
R7116 VDD.n297 VDD.n296 0.450111
R7117 VDD.n235 VDD.n234 0.449462
R7118 VDD.n354 VDD.n353 0.410734
R7119 VDD.n356 VDD.n355 0.410734
R7120 VDD.n440 VDD.n439 0.386525
R7121 VDD.n530 VDD.n505 0.359
R7122 VDD.n566 VDD.n530 0.359
R7123 VDD.n177 VDD.t174 0.3255
R7124 VDD.n177 VDD.t257 0.3255
R7125 VDD.n169 VDD.t214 0.3255
R7126 VDD.n169 VDD.t245 0.3255
R7127 VDD.n161 VDD.t157 0.3255
R7128 VDD.n161 VDD.t212 0.3255
R7129 VDD.n301 VDD.t180 0.3255
R7130 VDD.n301 VDD.t247 0.3255
R7131 VDD.n311 VDD.t259 0.3255
R7132 VDD.n311 VDD.t191 0.3255
R7133 VDD.n321 VDD.t249 0.3255
R7134 VDD.n321 VDD.t193 0.3255
R7135 VDD.n521 VDD.n520 0.305021
R7136 VDD.n367 VDD.n345 0.272055
R7137 VDD.n371 VDD.n340 0.272055
R7138 VDD.n372 VDD.n371 0.272055
R7139 VDD.n383 VDD.n375 0.272055
R7140 VDD.n522 VDD.n521 0.2705
R7141 VDD.n358 VDD.n357 0.242579
R7142 VDD.n258 VDD.n257 0.239643
R7143 VDD.n336 VDD.n335 0.21542
R7144 VDD.n440 VDD.n336 0.18923
R7145 VDD.n395 VDD.n394 0.181952
R7146 VDD.n7 VDD.n6 0.17077
R7147 VDD.n146 VDD.n7 0.17077
R7148 VDD.n105 VDD.n8 0.17077
R7149 VDD.n146 VDD.n8 0.17077
R7150 VDD.n343 VDD.n341 0.17077
R7151 VDD.n369 VDD.n343 0.17077
R7152 VDD.n344 VDD.n342 0.17077
R7153 VDD.n369 VDD.n342 0.17077
R7154 VDD.n378 VDD.n377 0.17077
R7155 VDD.n381 VDD.n377 0.17077
R7156 VDD.n376 VDD.n338 0.17077
R7157 VDD.n381 VDD.n376 0.17077
R7158 VDD.n552 VDD.n551 0.149678
R7159 VDD.n252 VDD.n251 0.149643
R7160 VDD.n251 VDD.n249 0.149643
R7161 VDD.n395 VDD.n393 0.146702
R7162 VDD.n519 VDD.n518 0.142281
R7163 VDD.n551 VDD.n550 0.131185
R7164 VDD.n253 VDD.n246 0.127143
R7165 VDD.n482 VDD.n481 0.126253
R7166 VDD.n523 VDD.n522 0.120089
R7167 VDD.n245 VDD.n244 0.120071
R7168 VDD.n365 VDD.n364 0.11975
R7169 VDD.n364 VDD.n363 0.11975
R7170 VDD.n363 VDD.n347 0.11975
R7171 VDD.n359 VDD.n347 0.11975
R7172 VDD.n366 VDD.n346 0.11975
R7173 VDD.n362 VDD.n346 0.11975
R7174 VDD.n362 VDD.n361 0.11975
R7175 VDD.n361 VDD.n360 0.11975
R7176 VDD.n390 VDD.n389 0.11975
R7177 VDD.n389 VDD.n388 0.11975
R7178 VDD.n388 VDD.n339 0.11975
R7179 VDD.n384 VDD.n339 0.11975
R7180 VDD.n391 VDD.n337 0.11975
R7181 VDD.n387 VDD.n337 0.11975
R7182 VDD.n387 VDD.n386 0.11975
R7183 VDD.n386 VDD.n385 0.11975
R7184 VDD.n480 VDD.n479 0.115158
R7185 VDD.n524 VDD.n523 0.113925
R7186 VDD.n554 VDD.n553 0.113925
R7187 VDD.n520 VDD.n519 0.10776
R7188 VDD.n36 VDD.n35 0.107449
R7189 VDD.n547 VDD.n546 0.106527
R7190 VDD.n184 VDD.n180 0.105016
R7191 VDD.n195 VDD.n180 0.105016
R7192 VDD.n197 VDD.n195 0.105016
R7193 VDD.n197 VDD.n196 0.105016
R7194 VDD.n196 VDD.n172 0.105016
R7195 VDD.n209 VDD.n172 0.105016
R7196 VDD.n211 VDD.n209 0.105016
R7197 VDD.n211 VDD.n210 0.105016
R7198 VDD.n210 VDD.n164 0.105016
R7199 VDD.n223 VDD.n164 0.105016
R7200 VDD.n226 VDD.n223 0.105016
R7201 VDD.n226 VDD.n225 0.105016
R7202 VDD.n225 VDD.n154 0.105016
R7203 VDD.n238 VDD.n154 0.105016
R7204 VDD.n496 VDD.n495 0.103753
R7205 VDD.n461 VDD.n460 0.101558
R7206 VDD.n549 VDD.n548 0.100363
R7207 VDD.n454 VDD.n453 0.0935717
R7208 VDD.n556 VDD.n555 0.0929658
R7209 VDD.n334 VDD.n333 0.0921268
R7210 VDD.n489 VDD.n488 0.0920411
R7211 VDD.n448 VDD.n447 0.0874283
R7212 VDD.n485 VDD.n484 0.080637
R7213 VDD.n95 VDD.n94 0.0794561
R7214 VDD.n450 VDD.n449 0.0791348
R7215 VDD.n559 VDD.n558 0.0757055
R7216 VDD.n446 VDD.n445 0.0751416
R7217 VDD.n558 VDD.n557 0.0744726
R7218 VDD.n498 VDD.n497 0.0723151
R7219 VDD.n493 VDD.n492 0.0692329
R7220 VDD.n336 VDD.n153 0.0672195
R7221 VDD.n458 VDD.n457 0.0671553
R7222 VDD.n555 VDD.n554 0.0646096
R7223 VDD.n445 VDD.n444 0.0634693
R7224 VDD.n525 VDD.n524 0.0624521
R7225 VDD.n561 VDD.n560 0.0624521
R7226 VDD.n452 VDD.n441 0.0622406
R7227 VDD.n367 VDD.n366 0.060125
R7228 VDD.n384 VDD.n383 0.060125
R7229 VDD.n385 VDD.n374 0.060125
R7230 VDD.n449 VDD.n448 0.0594761
R7231 VDD.n451 VDD.n450 0.0594761
R7232 VDD.n457 VDD.n456 0.0591689
R7233 VDD.n477 VDD.n476 0.0584452
R7234 VDD.n484 VDD.n483 0.0584452
R7235 VDD.n486 VDD.n485 0.0584452
R7236 VDD.n463 VDD.n451 0.0582474
R7237 VDD.n492 VDD.n491 0.0575205
R7238 VDD.n517 VDD.n516 0.0559795
R7239 VDD.n332 VDD.n278 0.0546935
R7240 VDD.n331 VDD.n263 0.0546935
R7241 VDD.n280 VDD.n277 0.0546935
R7242 VDD.n325 VDD.n264 0.0546935
R7243 VDD.n323 VDD.n276 0.0546935
R7244 VDD.n285 VDD.n265 0.0546935
R7245 VDD.n283 VDD.n275 0.0546935
R7246 VDD.n315 VDD.n266 0.0546935
R7247 VDD.n313 VDD.n274 0.0546935
R7248 VDD.n289 VDD.n267 0.0546935
R7249 VDD.n287 VDD.n273 0.0546935
R7250 VDD.n305 VDD.n268 0.0546935
R7251 VDD.n303 VDD.n272 0.0546935
R7252 VDD.n293 VDD.n269 0.0546935
R7253 VDD.n291 VDD.n271 0.0546935
R7254 VDD.n295 VDD.n270 0.0546935
R7255 VDD.n186 VDD.n185 0.0527581
R7256 VDD.n185 VDD.n183 0.0527581
R7257 VDD.n183 VDD.n181 0.0527581
R7258 VDD.n191 VDD.n181 0.0527581
R7259 VDD.n192 VDD.n191 0.0527581
R7260 VDD.n193 VDD.n192 0.0527581
R7261 VDD.n194 VDD.n193 0.0527581
R7262 VDD.n199 VDD.n198 0.0527581
R7263 VDD.n198 VDD.n179 0.0527581
R7264 VDD.n179 VDD.n173 0.0527581
R7265 VDD.n205 VDD.n173 0.0527581
R7266 VDD.n206 VDD.n205 0.0527581
R7267 VDD.n207 VDD.n206 0.0527581
R7268 VDD.n208 VDD.n207 0.0527581
R7269 VDD.n213 VDD.n212 0.0527581
R7270 VDD.n212 VDD.n171 0.0527581
R7271 VDD.n171 VDD.n165 0.0527581
R7272 VDD.n219 VDD.n165 0.0527581
R7273 VDD.n220 VDD.n219 0.0527581
R7274 VDD.n221 VDD.n220 0.0527581
R7275 VDD.n222 VDD.n221 0.0527581
R7276 VDD.n228 VDD.n227 0.0527581
R7277 VDD.n227 VDD.n163 0.0527581
R7278 VDD.n224 VDD.n163 0.0527581
R7279 VDD.n224 VDD.n158 0.0527581
R7280 VDD.n158 VDD.n157 0.0527581
R7281 VDD.n157 VDD.n155 0.0527581
R7282 VDD.n237 VDD.n155 0.0527581
R7283 VDD.n237 VDD.n236 0.0527581
R7284 VDD.n259 VDD.n245 0.0519286
R7285 VDD.n259 VDD.n258 0.0519286
R7286 VDD.n257 VDD.n256 0.0519286
R7287 VDD.n256 VDD.n246 0.0519286
R7288 VDD.n253 VDD.n252 0.0519286
R7289 VDD.n261 VDD.n240 0.0519286
R7290 VDD.n447 VDD.n446 0.0511826
R7291 VDD.n332 VDD.n331 0.0508226
R7292 VDD.n280 VDD.n263 0.0508226
R7293 VDD.n325 VDD.n277 0.0508226
R7294 VDD.n285 VDD.n276 0.0508226
R7295 VDD.n283 VDD.n265 0.0508226
R7296 VDD.n315 VDD.n275 0.0508226
R7297 VDD.n289 VDD.n274 0.0508226
R7298 VDD.n287 VDD.n267 0.0508226
R7299 VDD.n305 VDD.n273 0.0508226
R7300 VDD.n293 VDD.n272 0.0508226
R7301 VDD.n291 VDD.n269 0.0508226
R7302 VDD.n295 VDD.n271 0.0508226
R7303 VDD.n294 VDD.n270 0.0508226
R7304 VDD.n478 VDD.n477 0.0501233
R7305 VDD.n491 VDD.n490 0.0473493
R7306 VDD.n494 VDD.n493 0.0473493
R7307 VDD.n459 VDD.n458 0.0471894
R7308 VDD.n456 VDD.n455 0.0471894
R7309 VDD.n488 VDD.n487 0.0470411
R7310 VDD.n557 VDD.n556 0.0461164
R7311 VDD.n528 VDD.n527 0.0456716
R7312 VDD.n564 VDD.n563 0.0456716
R7313 VDD.n453 VDD.n452 0.0450393
R7314 VDD.n444 VDD.n443 0.0447321
R7315 VDD.n194 VDD.n178 0.0421129
R7316 VDD.n208 VDD.n170 0.0421129
R7317 VDD.n222 VDD.n162 0.0421129
R7318 VDD.n93 VDD.n92 0.04025
R7319 VDD.n92 VDD.n91 0.04025
R7320 VDD.n91 VDD.n12 0.04025
R7321 VDD.n87 VDD.n12 0.04025
R7322 VDD.n83 VDD.n15 0.04025
R7323 VDD.n79 VDD.n15 0.04025
R7324 VDD.n77 VDD.n76 0.04025
R7325 VDD.n76 VDD.n17 0.04025
R7326 VDD.n72 VDD.n17 0.04025
R7327 VDD.n70 VDD.n69 0.04025
R7328 VDD.n69 VDD.n20 0.04025
R7329 VDD.n65 VDD.n20 0.04025
R7330 VDD.n63 VDD.n62 0.04025
R7331 VDD.n62 VDD.n23 0.04025
R7332 VDD.n58 VDD.n23 0.04025
R7333 VDD.n58 VDD.n57 0.04025
R7334 VDD.n55 VDD.n26 0.04025
R7335 VDD.n51 VDD.n26 0.04025
R7336 VDD.n51 VDD.n50 0.04025
R7337 VDD.n48 VDD.n28 0.04025
R7338 VDD.n44 VDD.n43 0.04025
R7339 VDD.n43 VDD.n42 0.04025
R7340 VDD.n42 VDD.n32 0.04025
R7341 VDD.n38 VDD.n32 0.04025
R7342 VDD.n38 VDD.n37 0.04025
R7343 VDD.n94 VDD.n11 0.04025
R7344 VDD.n90 VDD.n11 0.04025
R7345 VDD.n90 VDD.n89 0.04025
R7346 VDD.n89 VDD.n88 0.04025
R7347 VDD.n88 VDD.n13 0.04025
R7348 VDD.n82 VDD.n13 0.04025
R7349 VDD.n82 VDD.n81 0.04025
R7350 VDD.n81 VDD.n80 0.04025
R7351 VDD.n80 VDD.n16 0.04025
R7352 VDD.n75 VDD.n16 0.04025
R7353 VDD.n75 VDD.n74 0.04025
R7354 VDD.n74 VDD.n73 0.04025
R7355 VDD.n73 VDD.n18 0.04025
R7356 VDD.n68 VDD.n18 0.04025
R7357 VDD.n68 VDD.n67 0.04025
R7358 VDD.n67 VDD.n66 0.04025
R7359 VDD.n66 VDD.n21 0.04025
R7360 VDD.n61 VDD.n21 0.04025
R7361 VDD.n61 VDD.n60 0.04025
R7362 VDD.n60 VDD.n59 0.04025
R7363 VDD.n59 VDD.n24 0.04025
R7364 VDD.n54 VDD.n24 0.04025
R7365 VDD.n54 VDD.n53 0.04025
R7366 VDD.n53 VDD.n52 0.04025
R7367 VDD.n52 VDD.n27 0.04025
R7368 VDD.n47 VDD.n27 0.04025
R7369 VDD.n47 VDD.n46 0.04025
R7370 VDD.n46 VDD.n45 0.04025
R7371 VDD.n45 VDD.n29 0.04025
R7372 VDD.n41 VDD.n29 0.04025
R7373 VDD.n41 VDD.n40 0.04025
R7374 VDD.n40 VDD.n39 0.04025
R7375 VDD.n39 VDD.n33 0.04025
R7376 VDD.n322 VDD.n264 0.0401774
R7377 VDD.n312 VDD.n266 0.0401774
R7378 VDD.n302 VDD.n268 0.0401774
R7379 VDD.n44 VDD.n31 0.039875
R7380 VDD.n548 VDD.n547 0.0387192
R7381 VDD.n560 VDD.n559 0.0387192
R7382 VDD.n56 VDD.n55 0.038375
R7383 VDD.n462 VDD.n461 0.0370529
R7384 VDD.n85 VDD.n84 0.035375
R7385 VDD.n497 VDD.n496 0.0353288
R7386 VDD.n490 VDD.n489 0.0347123
R7387 VDD.n86 VDD.n85 0.034625
R7388 VDD.n502 VDD.n500 0.0331712
R7389 VDD.n65 VDD.n64 0.033125
R7390 VDD.n455 VDD.n454 0.0327526
R7391 VDD.n546 VDD.n545 0.0325548
R7392 VDD.n499 VDD.n498 0.0322466
R7393 VDD.n526 VDD.n525 0.0322466
R7394 VDD.n562 VDD.n561 0.0322466
R7395 VDD.n465 VDD.n441 0.0321382
R7396 VDD.n466 VDD.n465 0.0318362
R7397 VDD.n143 VDD.n9 0.0306899
R7398 VDD.n139 VDD.n9 0.0306899
R7399 VDD.n139 VDD.n138 0.0306899
R7400 VDD.n138 VDD.n137 0.0306899
R7401 VDD.n137 VDD.n97 0.0306899
R7402 VDD.n133 VDD.n97 0.0306899
R7403 VDD.n133 VDD.n132 0.0306899
R7404 VDD.n132 VDD.n131 0.0306899
R7405 VDD.n131 VDD.n99 0.0306899
R7406 VDD.n127 VDD.n99 0.0306899
R7407 VDD.n127 VDD.n126 0.0306899
R7408 VDD.n126 VDD.n125 0.0306899
R7409 VDD.n125 VDD.n101 0.0306899
R7410 VDD.n121 VDD.n101 0.0306899
R7411 VDD.n121 VDD.n120 0.0306899
R7412 VDD.n120 VDD.n119 0.0306899
R7413 VDD.n119 VDD.n103 0.0306899
R7414 VDD.n115 VDD.n114 0.0306899
R7415 VDD.n114 VDD.n113 0.0306899
R7416 VDD.n113 VDD.n106 0.0306899
R7417 VDD.n109 VDD.n106 0.0306899
R7418 VDD.n109 VDD.n108 0.0306899
R7419 VDD.n108 VDD.n1 0.0306899
R7420 VDD.n583 VDD.n1 0.0306899
R7421 VDD.n583 VDD.n582 0.0306899
R7422 VDD.n582 VDD.n2 0.0306899
R7423 VDD.n578 VDD.n2 0.0306899
R7424 VDD.n578 VDD.n577 0.0306899
R7425 VDD.n577 VDD.n576 0.0306899
R7426 VDD.n576 VDD.n4 0.0306899
R7427 VDD.n572 VDD.n4 0.0306899
R7428 VDD.n572 VDD.n571 0.0306899
R7429 VDD.n571 VDD.n570 0.0306899
R7430 VDD.n570 VDD.n149 0.0306899
R7431 VDD.n49 VDD.n48 0.029375
R7432 VDD.n78 VDD.n77 0.025625
R7433 VDD.n553 VDD.n552 0.0251575
R7434 VDD.n460 VDD.n459 0.0247662
R7435 VDD.n72 VDD.n71 0.024125
R7436 VDD.n403 VDD.n402 0.024117
R7437 VDD.n410 VDD.n409 0.024117
R7438 VDD.n417 VDD.n416 0.024117
R7439 VDD.n424 VDD.n423 0.024117
R7440 VDD.n431 VDD.n430 0.024117
R7441 VDD.n438 VDD.n437 0.024117
R7442 VDD.n501 VDD.n469 0.0239247
R7443 VDD.n545 VDD.n544 0.0239247
R7444 VDD.n403 VDD.n398 0.0237979
R7445 VDD.n410 VDD.n405 0.0237979
R7446 VDD.n417 VDD.n412 0.0237979
R7447 VDD.n424 VDD.n419 0.0237979
R7448 VDD.n431 VDD.n426 0.0237979
R7449 VDD.n438 VDD.n433 0.0237979
R7450 VDD.n495 VDD.n494 0.023
R7451 VDD.n463 VDD.n462 0.0213874
R7452 VDD.n400 VDD.n399 0.020375
R7453 VDD.n401 VDD.n400 0.020375
R7454 VDD.n407 VDD.n406 0.020375
R7455 VDD.n408 VDD.n407 0.020375
R7456 VDD.n414 VDD.n413 0.020375
R7457 VDD.n415 VDD.n414 0.020375
R7458 VDD.n421 VDD.n420 0.020375
R7459 VDD.n422 VDD.n421 0.020375
R7460 VDD.n428 VDD.n427 0.020375
R7461 VDD.n429 VDD.n428 0.020375
R7462 VDD.n435 VDD.n434 0.020375
R7463 VDD.n436 VDD.n435 0.020375
R7464 VDD.n504 VDD.n468 0.0168356
R7465 VDD.n504 VDD.n503 0.0168356
R7466 VDD.n529 VDD.n506 0.0168356
R7467 VDD.n565 VDD.n531 0.0168356
R7468 VDD.n71 VDD.n70 0.016625
R7469 VDD.n105 VDD.n103 0.0161646
R7470 VDD.n79 VDD.n78 0.015125
R7471 VDD.n115 VDD.n105 0.0150253
R7472 VDD.n479 VDD.n478 0.0115959
R7473 VDD.n481 VDD.n480 0.0115959
R7474 VDD.n487 VDD.n486 0.0115959
R7475 VDD.n50 VDD.n49 0.011375
R7476 VDD.n199 VDD.n178 0.0111452
R7477 VDD.n213 VDD.n170 0.0111452
R7478 VDD.n228 VDD.n162 0.0111452
R7479 VDD.n323 VDD.n322 0.0111452
R7480 VDD.n313 VDD.n312 0.0111452
R7481 VDD.n303 VDD.n302 0.0111452
R7482 VDD.n483 VDD.n482 0.0100548
R7483 VDD.n142 VDD.n141 0.00804747
R7484 VDD.n141 VDD.n140 0.00804747
R7485 VDD.n140 VDD.n96 0.00804747
R7486 VDD.n136 VDD.n96 0.00804747
R7487 VDD.n136 VDD.n135 0.00804747
R7488 VDD.n135 VDD.n134 0.00804747
R7489 VDD.n134 VDD.n98 0.00804747
R7490 VDD.n130 VDD.n98 0.00804747
R7491 VDD.n130 VDD.n129 0.00804747
R7492 VDD.n129 VDD.n128 0.00804747
R7493 VDD.n128 VDD.n100 0.00804747
R7494 VDD.n124 VDD.n100 0.00804747
R7495 VDD.n124 VDD.n123 0.00804747
R7496 VDD.n123 VDD.n122 0.00804747
R7497 VDD.n122 VDD.n102 0.00804747
R7498 VDD.n118 VDD.n102 0.00804747
R7499 VDD.n118 VDD.n117 0.00804747
R7500 VDD.n117 VDD.n116 0.00804747
R7501 VDD.n116 VDD.n104 0.00804747
R7502 VDD.n112 VDD.n104 0.00804747
R7503 VDD.n112 VDD.n111 0.00804747
R7504 VDD.n111 VDD.n110 0.00804747
R7505 VDD.n110 VDD.n107 0.00804747
R7506 VDD.n107 VDD.n0 0.00804747
R7507 VDD.n584 VDD.n0 0.00804747
R7508 VDD.n581 VDD.n580 0.00804747
R7509 VDD.n580 VDD.n579 0.00804747
R7510 VDD.n579 VDD.n3 0.00804747
R7511 VDD.n575 VDD.n3 0.00804747
R7512 VDD.n575 VDD.n574 0.00804747
R7513 VDD.n574 VDD.n573 0.00804747
R7514 VDD.n573 VDD.n5 0.00804747
R7515 VDD.n569 VDD.n5 0.00804747
R7516 VDD.n569 VDD.n568 0.00804747
R7517 VDD.n550 VDD.n549 0.00789726
R7518 VDD.n64 VDD.n63 0.007625
R7519 VDD.n581 VDD 0.00754905
R7520 VDD.n87 VDD.n86 0.006125
R7521 VDD.n84 VDD.n83 0.005375
R7522 VDD.n248 VDD.n153 0.00522745
R7523 VDD.n248 VDD.n151 0.00522745
R7524 VDD.n262 VDD.n239 0.00481978
R7525 VDD.n239 VDD.n152 0.00481882
R7526 VDD.n93 VDD.n10 0.003875
R7527 VDD.n37 VDD.n36 0.003125
R7528 VDD.n518 VDD.n517 0.00296575
R7529 VDD.n57 VDD.n56 0.002375
R7530 VDD.n500 VDD.n499 0.00142466
R7531 VDD.n502 VDD.n501 0.00142466
R7532 VDD.n527 VDD.n526 0.00142466
R7533 VDD.n563 VDD.n562 0.00142466
R7534 VDD.n584 VDD 0.000998418
R7535 VDD.n31 VDD.n28 0.000875
R7536 a_24355_n1338.n0 a_24355_n1338.t41 14.4185
R7537 a_24355_n1338.n1 a_24355_n1338.t50 14.4185
R7538 a_24355_n1338.n0 a_24355_n1338.n23 11.7725
R7539 a_24355_n1338.n0 a_24355_n1338.n21 11.7725
R7540 a_24355_n1338.n0 a_24355_n1338.n19 11.7725
R7541 a_24355_n1338.n0 a_24355_n1338.n17 11.7725
R7542 a_24355_n1338.n0 a_24355_n1338.n15 11.7725
R7543 a_24355_n1338.n1 a_24355_n1338.n13 11.7725
R7544 a_24355_n1338.n1 a_24355_n1338.n11 11.7725
R7545 a_24355_n1338.n1 a_24355_n1338.n9 11.7725
R7546 a_24355_n1338.n1 a_24355_n1338.n7 11.7725
R7547 a_24355_n1338.n3 a_24355_n1338.n26 7.13263
R7548 a_24355_n1338.n3 a_24355_n1338.n4 6.43746
R7549 a_24355_n1338.n3 a_24355_n1338.n25 6.43746
R7550 a_24355_n1338.n3 a_24355_n1338.n6 6.43746
R7551 a_24355_n1338.n0 a_24355_n1338.t44 3.93079
R7552 a_24355_n1338.n1 a_24355_n1338.t15 3.93079
R7553 a_24355_n1338.n4 a_24355_n1338.t26 3.8098
R7554 a_24355_n1338.n4 a_24355_n1338.t20 3.8098
R7555 a_24355_n1338.n26 a_24355_n1338.t21 3.8098
R7556 a_24355_n1338.n26 a_24355_n1338.t22 3.8098
R7557 a_24355_n1338.n25 a_24355_n1338.t25 3.8098
R7558 a_24355_n1338.n25 a_24355_n1338.t27 3.8098
R7559 a_24355_n1338.n6 a_24355_n1338.t23 3.8098
R7560 a_24355_n1338.n6 a_24355_n1338.t24 3.8098
R7561 a_24355_n1338.n2 a_24355_n1338.n28 3.34593
R7562 a_24355_n1338.n0 a_24355_n1338.n24 2.95079
R7563 a_24355_n1338.n0 a_24355_n1338.n22 2.95079
R7564 a_24355_n1338.n0 a_24355_n1338.n20 2.95079
R7565 a_24355_n1338.n0 a_24355_n1338.n18 2.95079
R7566 a_24355_n1338.n0 a_24355_n1338.n16 2.95079
R7567 a_24355_n1338.n1 a_24355_n1338.n14 2.95079
R7568 a_24355_n1338.n1 a_24355_n1338.n12 2.95079
R7569 a_24355_n1338.n1 a_24355_n1338.n10 2.95079
R7570 a_24355_n1338.n1 a_24355_n1338.n8 2.95079
R7571 a_24355_n1338.n2 a_24355_n1338.n27 2.71593
R7572 a_24355_n1338.n3 a_24355_n1338.n5 2.71593
R7573 a_24355_n1338.n29 a_24355_n1338.n3 2.71593
R7574 a_24355_n1338.n27 a_24355_n1338.t28 2.06607
R7575 a_24355_n1338.n27 a_24355_n1338.t33 2.06607
R7576 a_24355_n1338.n28 a_24355_n1338.t31 2.06607
R7577 a_24355_n1338.n28 a_24355_n1338.t29 2.06607
R7578 a_24355_n1338.n5 a_24355_n1338.t34 2.06607
R7579 a_24355_n1338.n5 a_24355_n1338.t32 2.06607
R7580 a_24355_n1338.n29 a_24355_n1338.t30 2.06607
R7581 a_24355_n1338.t35 a_24355_n1338.n29 2.06607
R7582 a_24355_n1338.n23 a_24355_n1338.t13 1.6385
R7583 a_24355_n1338.n23 a_24355_n1338.t37 1.6385
R7584 a_24355_n1338.n21 a_24355_n1338.t42 1.6385
R7585 a_24355_n1338.n21 a_24355_n1338.t6 1.6385
R7586 a_24355_n1338.n19 a_24355_n1338.t19 1.6385
R7587 a_24355_n1338.n19 a_24355_n1338.t51 1.6385
R7588 a_24355_n1338.n17 a_24355_n1338.t18 1.6385
R7589 a_24355_n1338.n17 a_24355_n1338.t17 1.6385
R7590 a_24355_n1338.n15 a_24355_n1338.t3 1.6385
R7591 a_24355_n1338.n15 a_24355_n1338.t4 1.6385
R7592 a_24355_n1338.n13 a_24355_n1338.t11 1.6385
R7593 a_24355_n1338.n13 a_24355_n1338.t36 1.6385
R7594 a_24355_n1338.n11 a_24355_n1338.t5 1.6385
R7595 a_24355_n1338.n11 a_24355_n1338.t12 1.6385
R7596 a_24355_n1338.n9 a_24355_n1338.t38 1.6385
R7597 a_24355_n1338.n9 a_24355_n1338.t43 1.6385
R7598 a_24355_n1338.n7 a_24355_n1338.t7 1.6385
R7599 a_24355_n1338.n7 a_24355_n1338.t49 1.6385
R7600 a_24355_n1338.n3 a_24355_n1338.n1 1.61746
R7601 a_24355_n1338.n1 a_24355_n1338.n0 1.5593
R7602 a_24355_n1338.n3 a_24355_n1338.n2 0.925734
R7603 a_24355_n1338.n24 a_24355_n1338.t14 0.607167
R7604 a_24355_n1338.n24 a_24355_n1338.t45 0.607167
R7605 a_24355_n1338.n22 a_24355_n1338.t10 0.607167
R7606 a_24355_n1338.n22 a_24355_n1338.t39 0.607167
R7607 a_24355_n1338.n20 a_24355_n1338.t47 0.607167
R7608 a_24355_n1338.n20 a_24355_n1338.t2 0.607167
R7609 a_24355_n1338.n18 a_24355_n1338.t1 0.607167
R7610 a_24355_n1338.n18 a_24355_n1338.t55 0.607167
R7611 a_24355_n1338.n16 a_24355_n1338.t48 0.607167
R7612 a_24355_n1338.n16 a_24355_n1338.t16 0.607167
R7613 a_24355_n1338.n14 a_24355_n1338.t9 0.607167
R7614 a_24355_n1338.n14 a_24355_n1338.t53 0.607167
R7615 a_24355_n1338.n12 a_24355_n1338.t52 0.607167
R7616 a_24355_n1338.n12 a_24355_n1338.t0 0.607167
R7617 a_24355_n1338.n10 a_24355_n1338.t54 0.607167
R7618 a_24355_n1338.n10 a_24355_n1338.t46 0.607167
R7619 a_24355_n1338.n8 a_24355_n1338.t40 0.607167
R7620 a_24355_n1338.n8 a_24355_n1338.t8 0.607167
R7621 a_27899_438.t29 a_27899_438.n27 36.5005
R7622 a_27899_438.n10 a_27899_438.t16 36.5005
R7623 a_27899_438.n28 a_27899_438.t29 33.21
R7624 a_27899_438.t16 a_27899_438.n9 33.21
R7625 a_27899_438.n11 a_27899_438.n10 18.8035
R7626 a_27899_438.n12 a_27899_438.n11 18.8035
R7627 a_27899_438.n13 a_27899_438.n12 18.8035
R7628 a_27899_438.n14 a_27899_438.n13 18.8035
R7629 a_27899_438.n15 a_27899_438.n14 18.8035
R7630 a_27899_438.n16 a_27899_438.n15 18.8035
R7631 a_27899_438.n17 a_27899_438.n16 18.8035
R7632 a_27899_438.n18 a_27899_438.n17 18.8035
R7633 a_27899_438.n19 a_27899_438.n18 18.8035
R7634 a_27899_438.n20 a_27899_438.n19 18.8035
R7635 a_27899_438.n21 a_27899_438.n20 18.8035
R7636 a_27899_438.n22 a_27899_438.n21 18.8035
R7637 a_27899_438.n23 a_27899_438.n22 18.8035
R7638 a_27899_438.n24 a_27899_438.n23 18.8035
R7639 a_27899_438.n25 a_27899_438.n24 18.8035
R7640 a_27899_438.n26 a_27899_438.n25 18.8035
R7641 a_27899_438.n27 a_27899_438.n26 18.8035
R7642 a_27899_438.n9 a_27899_438.t21 17.6975
R7643 a_27899_438.n10 a_27899_438.t21 17.6975
R7644 a_27899_438.n8 a_27899_438.t14 17.6975
R7645 a_27899_438.n11 a_27899_438.t14 17.6975
R7646 a_27899_438.n7 a_27899_438.t17 17.6975
R7647 a_27899_438.n12 a_27899_438.t17 17.6975
R7648 a_27899_438.n6 a_27899_438.t31 17.6975
R7649 a_27899_438.n13 a_27899_438.t31 17.6975
R7650 a_27899_438.n5 a_27899_438.t27 17.6975
R7651 a_27899_438.n14 a_27899_438.t27 17.6975
R7652 a_27899_438.n4 a_27899_438.t30 17.6975
R7653 a_27899_438.n15 a_27899_438.t30 17.6975
R7654 a_27899_438.n3 a_27899_438.t26 17.6975
R7655 a_27899_438.n16 a_27899_438.t26 17.6975
R7656 a_27899_438.n2 a_27899_438.t25 17.6975
R7657 a_27899_438.n17 a_27899_438.t25 17.6975
R7658 a_27899_438.t22 a_27899_438.n1 17.6975
R7659 a_27899_438.n18 a_27899_438.t22 17.6975
R7660 a_27899_438.n36 a_27899_438.t23 17.6975
R7661 a_27899_438.n19 a_27899_438.t23 17.6975
R7662 a_27899_438.n35 a_27899_438.t19 17.6975
R7663 a_27899_438.n20 a_27899_438.t19 17.6975
R7664 a_27899_438.n34 a_27899_438.t13 17.6975
R7665 a_27899_438.n21 a_27899_438.t13 17.6975
R7666 a_27899_438.n33 a_27899_438.t24 17.6975
R7667 a_27899_438.n22 a_27899_438.t24 17.6975
R7668 a_27899_438.n32 a_27899_438.t20 17.6975
R7669 a_27899_438.n23 a_27899_438.t20 17.6975
R7670 a_27899_438.n31 a_27899_438.t15 17.6975
R7671 a_27899_438.n24 a_27899_438.t15 17.6975
R7672 a_27899_438.n30 a_27899_438.t18 17.6975
R7673 a_27899_438.n25 a_27899_438.t18 17.6975
R7674 a_27899_438.n29 a_27899_438.t32 17.6975
R7675 a_27899_438.n26 a_27899_438.t32 17.6975
R7676 a_27899_438.n28 a_27899_438.t28 17.6975
R7677 a_27899_438.n27 a_27899_438.t28 17.6975
R7678 a_27899_438.n9 a_27899_438.n8 15.513
R7679 a_27899_438.n8 a_27899_438.n7 15.513
R7680 a_27899_438.n7 a_27899_438.n6 15.513
R7681 a_27899_438.n6 a_27899_438.n5 15.513
R7682 a_27899_438.n5 a_27899_438.n4 15.513
R7683 a_27899_438.n4 a_27899_438.n3 15.513
R7684 a_27899_438.n3 a_27899_438.n2 15.513
R7685 a_27899_438.n2 a_27899_438.n1 15.513
R7686 a_27899_438.n36 a_27899_438.n35 15.513
R7687 a_27899_438.n35 a_27899_438.n34 15.513
R7688 a_27899_438.n34 a_27899_438.n33 15.513
R7689 a_27899_438.n33 a_27899_438.n32 15.513
R7690 a_27899_438.n32 a_27899_438.n31 15.513
R7691 a_27899_438.n31 a_27899_438.n30 15.513
R7692 a_27899_438.n30 a_27899_438.n29 15.513
R7693 a_27899_438.n29 a_27899_438.n28 15.513
R7694 a_27899_438.n0 a_27899_438.n1 7.75675
R7695 a_27899_438.n0 a_27899_438.n36 7.75675
R7696 a_27899_438.n0 a_27899_438.t7 6.85374
R7697 a_27899_438.n0 a_27899_438.t6 6.41398
R7698 a_27899_438.n0 a_27899_438.t0 6.41398
R7699 a_27899_438.n0 a_27899_438.t5 5.44249
R7700 a_27899_438.n0 a_27899_438.t10 4.78346
R7701 a_27899_438.n0 a_27899_438.t9 4.78151
R7702 a_27899_438.t1 a_27899_438.n37 2.06607
R7703 a_27899_438.n37 a_27899_438.t12 2.06607
R7704 a_27899_438.t6 a_27899_438.t2 1.99806
R7705 a_27899_438.t7 a_27899_438.t11 1.99806
R7706 a_27899_438.t3 a_27899_438.t4 1.99806
R7707 a_27899_438.t0 a_27899_438.t8 1.99806
R7708 a_27899_438.n0 a_27899_438.t3 7.1833
R7709 a_27899_438.n37 a_27899_438.n0 5.56319
R7710 PLL_CLK_OUT.n11 PLL_CLK_OUT.n10 15.3005
R7711 PLL_CLK_OUT.n13 PLL_CLK_OUT.n12 15.3005
R7712 PLL_CLK_OUT.n15 PLL_CLK_OUT.n14 15.3005
R7713 PLL_CLK_OUT.n17 PLL_CLK_OUT.n16 15.3005
R7714 PLL_CLK_OUT.n19 PLL_CLK_OUT.n18 15.3005
R7715 PLL_CLK_OUT.n21 PLL_CLK_OUT.n20 15.3005
R7716 PLL_CLK_OUT.n23 PLL_CLK_OUT.n22 15.3005
R7717 PLL_CLK_OUT.n25 PLL_CLK_OUT.n24 15.3005
R7718 PLL_CLK_OUT.n27 PLL_CLK_OUT.n26 15.3005
R7719 PLL_CLK_OUT.n29 PLL_CLK_OUT.n28 15.3005
R7720 PLL_CLK_OUT.n11 PLL_CLK_OUT.n9 5.21417
R7721 PLL_CLK_OUT.n13 PLL_CLK_OUT.n8 5.21417
R7722 PLL_CLK_OUT.n15 PLL_CLK_OUT.n7 5.21417
R7723 PLL_CLK_OUT.n17 PLL_CLK_OUT.n6 5.21417
R7724 PLL_CLK_OUT.n19 PLL_CLK_OUT.n5 5.21417
R7725 PLL_CLK_OUT.n21 PLL_CLK_OUT.n4 5.21417
R7726 PLL_CLK_OUT.n23 PLL_CLK_OUT.n3 5.21417
R7727 PLL_CLK_OUT.n25 PLL_CLK_OUT.n2 5.21417
R7728 PLL_CLK_OUT.n27 PLL_CLK_OUT.n1 5.21417
R7729 PLL_CLK_OUT.n29 PLL_CLK_OUT.n0 5.21417
R7730 PLL_CLK_OUT PLL_CLK_OUT.n29 1.71725
R7731 PLL_CLK_OUT.n10 PLL_CLK_OUT.t13 1.6385
R7732 PLL_CLK_OUT.n10 PLL_CLK_OUT.t12 1.6385
R7733 PLL_CLK_OUT.n12 PLL_CLK_OUT.t23 1.6385
R7734 PLL_CLK_OUT.n12 PLL_CLK_OUT.t9 1.6385
R7735 PLL_CLK_OUT.n14 PLL_CLK_OUT.t21 1.6385
R7736 PLL_CLK_OUT.n14 PLL_CLK_OUT.t26 1.6385
R7737 PLL_CLK_OUT.n16 PLL_CLK_OUT.t28 1.6385
R7738 PLL_CLK_OUT.n16 PLL_CLK_OUT.t17 1.6385
R7739 PLL_CLK_OUT.n18 PLL_CLK_OUT.t18 1.6385
R7740 PLL_CLK_OUT.n18 PLL_CLK_OUT.t22 1.6385
R7741 PLL_CLK_OUT.n20 PLL_CLK_OUT.t16 1.6385
R7742 PLL_CLK_OUT.n20 PLL_CLK_OUT.t19 1.6385
R7743 PLL_CLK_OUT.n22 PLL_CLK_OUT.t11 1.6385
R7744 PLL_CLK_OUT.n22 PLL_CLK_OUT.t15 1.6385
R7745 PLL_CLK_OUT.n24 PLL_CLK_OUT.t10 1.6385
R7746 PLL_CLK_OUT.n24 PLL_CLK_OUT.t14 1.6385
R7747 PLL_CLK_OUT.n26 PLL_CLK_OUT.t27 1.6385
R7748 PLL_CLK_OUT.n26 PLL_CLK_OUT.t24 1.6385
R7749 PLL_CLK_OUT.n28 PLL_CLK_OUT.t25 1.6385
R7750 PLL_CLK_OUT.n28 PLL_CLK_OUT.t20 1.6385
R7751 PLL_CLK_OUT.n9 PLL_CLK_OUT.t3 0.607167
R7752 PLL_CLK_OUT.n9 PLL_CLK_OUT.t7 0.607167
R7753 PLL_CLK_OUT.n8 PLL_CLK_OUT.t33 0.607167
R7754 PLL_CLK_OUT.n8 PLL_CLK_OUT.t30 0.607167
R7755 PLL_CLK_OUT.n7 PLL_CLK_OUT.t0 0.607167
R7756 PLL_CLK_OUT.n7 PLL_CLK_OUT.t38 0.607167
R7757 PLL_CLK_OUT.n6 PLL_CLK_OUT.t37 0.607167
R7758 PLL_CLK_OUT.n6 PLL_CLK_OUT.t36 0.607167
R7759 PLL_CLK_OUT.n5 PLL_CLK_OUT.t8 0.607167
R7760 PLL_CLK_OUT.n5 PLL_CLK_OUT.t4 0.607167
R7761 PLL_CLK_OUT.n4 PLL_CLK_OUT.t39 0.607167
R7762 PLL_CLK_OUT.n4 PLL_CLK_OUT.t35 0.607167
R7763 PLL_CLK_OUT.n3 PLL_CLK_OUT.t2 0.607167
R7764 PLL_CLK_OUT.n3 PLL_CLK_OUT.t1 0.607167
R7765 PLL_CLK_OUT.n2 PLL_CLK_OUT.t29 0.607167
R7766 PLL_CLK_OUT.n2 PLL_CLK_OUT.t34 0.607167
R7767 PLL_CLK_OUT.n1 PLL_CLK_OUT.t32 0.607167
R7768 PLL_CLK_OUT.n1 PLL_CLK_OUT.t5 0.607167
R7769 PLL_CLK_OUT.n0 PLL_CLK_OUT.t31 0.607167
R7770 PLL_CLK_OUT.n0 PLL_CLK_OUT.t6 0.607167
R7771 PLL_CLK_OUT.n29 PLL_CLK_OUT.n27 0.1535
R7772 PLL_CLK_OUT.n27 PLL_CLK_OUT.n25 0.1535
R7773 PLL_CLK_OUT.n25 PLL_CLK_OUT.n23 0.1535
R7774 PLL_CLK_OUT.n23 PLL_CLK_OUT.n21 0.1535
R7775 PLL_CLK_OUT.n21 PLL_CLK_OUT.n19 0.1535
R7776 PLL_CLK_OUT.n19 PLL_CLK_OUT.n17 0.1535
R7777 PLL_CLK_OUT.n17 PLL_CLK_OUT.n15 0.1535
R7778 PLL_CLK_OUT.n15 PLL_CLK_OUT.n13 0.1535
R7779 PLL_CLK_OUT.n13 PLL_CLK_OUT.n11 0.1535
R7780 a_5840_15093.t9 a_5840_15093.t4 29.4935
R7781 a_5840_15093.n35 a_5840_15093.n112 11.0705
R7782 a_5840_15093.n35 a_5840_15093.n111 11.0705
R7783 a_5840_15093.n34 a_5840_15093.n37 1.49211
R7784 a_5840_15093.n36 a_5840_15093.n34 2.24415
R7785 a_5840_15093.n35 a_5840_15093.n39 2.24276
R7786 a_5840_15093.n36 a_5840_15093.n39 0.0174769
R7787 a_5840_15093.n34 a_5840_15093.n41 4.27695
R7788 a_5840_15093.n113 a_5840_15093.n34 4.27695
R7789 a_5840_15093.n40 a_5840_15093.n37 0.0102449
R7790 a_5840_15093.n35 a_5840_15093.n38 2.24438
R7791 a_5840_15093.n112 a_5840_15093.t7 1.6385
R7792 a_5840_15093.n112 a_5840_15093.t6 1.6385
R7793 a_5840_15093.n111 a_5840_15093.t8 1.6385
R7794 a_5840_15093.n111 a_5840_15093.t5 1.6385
R7795 a_5840_15093.n3 a_5840_15093.n36 1.51491
R7796 a_5840_15093.n108 a_5840_15093.n0 1.5005
R7797 a_5840_15093.n107 a_5840_15093.n6 0.0148215
R7798 a_5840_15093.n0 a_5840_15093.n6 0.744089
R7799 a_5840_15093.n103 a_5840_15093.n7 0.0148215
R7800 a_5840_15093.n7 a_5840_15093.n0 0.744089
R7801 a_5840_15093.n101 a_5840_15093.n9 0.0148215
R7802 a_5840_15093.n0 a_5840_15093.n9 0.744089
R7803 a_5840_15093.n97 a_5840_15093.n10 0.0148215
R7804 a_5840_15093.n10 a_5840_15093.n0 0.744089
R7805 a_5840_15093.n95 a_5840_15093.n12 0.0148215
R7806 a_5840_15093.n0 a_5840_15093.n12 0.744089
R7807 a_5840_15093.n91 a_5840_15093.n13 0.0148215
R7808 a_5840_15093.n13 a_5840_15093.n0 0.744089
R7809 a_5840_15093.n89 a_5840_15093.n15 0.0148215
R7810 a_5840_15093.n0 a_5840_15093.n15 0.744089
R7811 a_5840_15093.n85 a_5840_15093.n16 0.0148215
R7812 a_5840_15093.n16 a_5840_15093.n0 0.744089
R7813 a_5840_15093.n83 a_5840_15093.n18 0.0148215
R7814 a_5840_15093.n0 a_5840_15093.n18 0.744089
R7815 a_5840_15093.n79 a_5840_15093.n19 0.0148215
R7816 a_5840_15093.n19 a_5840_15093.n0 0.744089
R7817 a_5840_15093.n77 a_5840_15093.n21 0.0148215
R7818 a_5840_15093.n0 a_5840_15093.n21 0.744089
R7819 a_5840_15093.n73 a_5840_15093.n22 0.0148215
R7820 a_5840_15093.n22 a_5840_15093.n1 0.744089
R7821 a_5840_15093.n71 a_5840_15093.n24 0.0148215
R7822 a_5840_15093.n1 a_5840_15093.n24 0.744089
R7823 a_5840_15093.n67 a_5840_15093.n25 0.0148215
R7824 a_5840_15093.n25 a_5840_15093.n1 0.744089
R7825 a_5840_15093.n65 a_5840_15093.n27 0.0148215
R7826 a_5840_15093.n1 a_5840_15093.n27 0.744089
R7827 a_5840_15093.n61 a_5840_15093.n28 0.0148215
R7828 a_5840_15093.n28 a_5840_15093.n1 0.744089
R7829 a_5840_15093.n59 a_5840_15093.n30 0.0148215
R7830 a_5840_15093.n1 a_5840_15093.n30 0.744089
R7831 a_5840_15093.n55 a_5840_15093.n31 0.0148215
R7832 a_5840_15093.n31 a_5840_15093.n1 0.744089
R7833 a_5840_15093.n53 a_5840_15093.n32 0.0148215
R7834 a_5840_15093.n1 a_5840_15093.n32 0.744089
R7835 a_5840_15093.n40 a_5840_15093.n3 1.5005
R7836 a_5840_15093.n3 a_5840_15093.n33 0.744089
R7837 a_5840_15093.n110 a_5840_15093.n109 1.5005
R7838 a_5840_15093.n108 a_5840_15093.n42 1.5005
R7839 a_5840_15093.n107 a_5840_15093.n106 1.5005
R7840 a_5840_15093.n105 a_5840_15093.n5 1.5005
R7841 a_5840_15093.n104 a_5840_15093.n103 1.5005
R7842 a_5840_15093.n102 a_5840_15093.n43 1.5005
R7843 a_5840_15093.n101 a_5840_15093.n100 1.5005
R7844 a_5840_15093.n99 a_5840_15093.n8 1.5005
R7845 a_5840_15093.n98 a_5840_15093.n97 1.5005
R7846 a_5840_15093.n96 a_5840_15093.n44 1.5005
R7847 a_5840_15093.n95 a_5840_15093.n94 1.5005
R7848 a_5840_15093.n93 a_5840_15093.n11 1.5005
R7849 a_5840_15093.n92 a_5840_15093.n91 1.5005
R7850 a_5840_15093.n90 a_5840_15093.n45 1.5005
R7851 a_5840_15093.n89 a_5840_15093.n88 1.5005
R7852 a_5840_15093.n87 a_5840_15093.n14 1.5005
R7853 a_5840_15093.n86 a_5840_15093.n85 1.5005
R7854 a_5840_15093.n84 a_5840_15093.n46 1.5005
R7855 a_5840_15093.n83 a_5840_15093.n82 1.5005
R7856 a_5840_15093.n81 a_5840_15093.n17 1.5005
R7857 a_5840_15093.n80 a_5840_15093.n79 1.5005
R7858 a_5840_15093.n78 a_5840_15093.n47 1.5005
R7859 a_5840_15093.n77 a_5840_15093.n76 1.5005
R7860 a_5840_15093.n75 a_5840_15093.n20 1.5005
R7861 a_5840_15093.n74 a_5840_15093.n73 1.5005
R7862 a_5840_15093.n72 a_5840_15093.n48 1.5005
R7863 a_5840_15093.n71 a_5840_15093.n70 1.5005
R7864 a_5840_15093.n69 a_5840_15093.n23 1.5005
R7865 a_5840_15093.n68 a_5840_15093.n67 1.5005
R7866 a_5840_15093.n66 a_5840_15093.n49 1.5005
R7867 a_5840_15093.n65 a_5840_15093.n64 1.5005
R7868 a_5840_15093.n63 a_5840_15093.n26 1.5005
R7869 a_5840_15093.n62 a_5840_15093.n61 1.5005
R7870 a_5840_15093.n60 a_5840_15093.n50 1.5005
R7871 a_5840_15093.n59 a_5840_15093.n58 1.5005
R7872 a_5840_15093.n57 a_5840_15093.n29 1.5005
R7873 a_5840_15093.n56 a_5840_15093.n55 1.5005
R7874 a_5840_15093.n54 a_5840_15093.n51 1.5005
R7875 a_5840_15093.n53 a_5840_15093.n52 1.5005
R7876 a_5840_15093.n41 a_5840_15093.t0 0.9105
R7877 a_5840_15093.n41 a_5840_15093.t1 0.9105
R7878 a_5840_15093.t3 a_5840_15093.n113 0.9105
R7879 a_5840_15093.n113 a_5840_15093.t2 0.9105
R7880 a_5840_15093.n1 a_5840_15093.n0 0.5213
R7881 a_5840_15093.n40 a_5840_15093.n39 0.0174769
R7882 a_5840_15093.n37 a_5840_15093.n38 0.0195402
R7883 a_5840_15093.n109 a_5840_15093.n108 0.0284
R7884 a_5840_15093.n108 a_5840_15093.n107 0.0284
R7885 a_5840_15093.n6 a_5840_15093.n5 0.0148215
R7886 a_5840_15093.n103 a_5840_15093.n5 0.0284
R7887 a_5840_15093.n7 a_5840_15093.n102 0.0148215
R7888 a_5840_15093.n102 a_5840_15093.n101 0.0284
R7889 a_5840_15093.n9 a_5840_15093.n8 0.0148215
R7890 a_5840_15093.n97 a_5840_15093.n8 0.0284
R7891 a_5840_15093.n10 a_5840_15093.n96 0.0148215
R7892 a_5840_15093.n96 a_5840_15093.n95 0.0284
R7893 a_5840_15093.n12 a_5840_15093.n11 0.0148215
R7894 a_5840_15093.n91 a_5840_15093.n11 0.0284
R7895 a_5840_15093.n13 a_5840_15093.n90 0.0148215
R7896 a_5840_15093.n90 a_5840_15093.n89 0.0284
R7897 a_5840_15093.n15 a_5840_15093.n14 0.0148215
R7898 a_5840_15093.n85 a_5840_15093.n14 0.0284
R7899 a_5840_15093.n16 a_5840_15093.n84 0.0148215
R7900 a_5840_15093.n84 a_5840_15093.n83 0.0284
R7901 a_5840_15093.n18 a_5840_15093.n17 0.0148215
R7902 a_5840_15093.n79 a_5840_15093.n17 0.0284
R7903 a_5840_15093.n19 a_5840_15093.n78 0.0148215
R7904 a_5840_15093.n78 a_5840_15093.n77 0.0284
R7905 a_5840_15093.n21 a_5840_15093.n20 0.0148215
R7906 a_5840_15093.n73 a_5840_15093.n20 0.0284
R7907 a_5840_15093.n22 a_5840_15093.n72 0.0148215
R7908 a_5840_15093.n72 a_5840_15093.n71 0.0284
R7909 a_5840_15093.n24 a_5840_15093.n23 0.0148215
R7910 a_5840_15093.n67 a_5840_15093.n23 0.0284
R7911 a_5840_15093.n25 a_5840_15093.n66 0.0148215
R7912 a_5840_15093.n66 a_5840_15093.n65 0.0284
R7913 a_5840_15093.n27 a_5840_15093.n26 0.0148215
R7914 a_5840_15093.n61 a_5840_15093.n26 0.0284
R7915 a_5840_15093.n28 a_5840_15093.n60 0.0148215
R7916 a_5840_15093.n60 a_5840_15093.n59 0.0284
R7917 a_5840_15093.n30 a_5840_15093.n29 0.0148215
R7918 a_5840_15093.n55 a_5840_15093.n29 0.0284
R7919 a_5840_15093.n31 a_5840_15093.n54 0.0148215
R7920 a_5840_15093.n54 a_5840_15093.n53 0.0284
R7921 a_5840_15093.n32 a_5840_15093.n2 0.0830103
R7922 a_5840_15093.n38 a_5840_15093.n33 0.0148215
R7923 a_5840_15093.n33 a_5840_15093.n110 0.0427215
R7924 a_5840_15093.n110 a_5840_15093.n42 0.0284
R7925 a_5840_15093.n106 a_5840_15093.n42 0.0284
R7926 a_5840_15093.n106 a_5840_15093.n105 0.0284
R7927 a_5840_15093.n105 a_5840_15093.n104 0.0284
R7928 a_5840_15093.n104 a_5840_15093.n43 0.0284
R7929 a_5840_15093.n100 a_5840_15093.n43 0.0284
R7930 a_5840_15093.n100 a_5840_15093.n99 0.0284
R7931 a_5840_15093.n99 a_5840_15093.n98 0.0284
R7932 a_5840_15093.n98 a_5840_15093.n44 0.0284
R7933 a_5840_15093.n94 a_5840_15093.n44 0.0284
R7934 a_5840_15093.n94 a_5840_15093.n93 0.0284
R7935 a_5840_15093.n93 a_5840_15093.n92 0.0284
R7936 a_5840_15093.n92 a_5840_15093.n45 0.0284
R7937 a_5840_15093.n88 a_5840_15093.n45 0.0284
R7938 a_5840_15093.n88 a_5840_15093.n87 0.0284
R7939 a_5840_15093.n87 a_5840_15093.n86 0.0284
R7940 a_5840_15093.n86 a_5840_15093.n46 0.0284
R7941 a_5840_15093.n82 a_5840_15093.n46 0.0284
R7942 a_5840_15093.n82 a_5840_15093.n81 0.0284
R7943 a_5840_15093.n81 a_5840_15093.n80 0.0284
R7944 a_5840_15093.n80 a_5840_15093.n47 0.0284
R7945 a_5840_15093.n76 a_5840_15093.n47 0.0284
R7946 a_5840_15093.n76 a_5840_15093.n75 0.0284
R7947 a_5840_15093.n75 a_5840_15093.n74 0.0284
R7948 a_5840_15093.n74 a_5840_15093.n48 0.0284
R7949 a_5840_15093.n70 a_5840_15093.n48 0.0284
R7950 a_5840_15093.n70 a_5840_15093.n69 0.0284
R7951 a_5840_15093.n69 a_5840_15093.n68 0.0284
R7952 a_5840_15093.n68 a_5840_15093.n49 0.0284
R7953 a_5840_15093.n64 a_5840_15093.n49 0.0284
R7954 a_5840_15093.n64 a_5840_15093.n63 0.0284
R7955 a_5840_15093.n63 a_5840_15093.n62 0.0284
R7956 a_5840_15093.n62 a_5840_15093.n50 0.0284
R7957 a_5840_15093.n58 a_5840_15093.n50 0.0284
R7958 a_5840_15093.n58 a_5840_15093.n57 0.0284
R7959 a_5840_15093.n57 a_5840_15093.n56 0.0284
R7960 a_5840_15093.n56 a_5840_15093.n51 0.0284
R7961 a_5840_15093.n52 a_5840_15093.n51 0.0284
R7962 a_5840_15093.n52 a_5840_15093.n2 0.23658
R7963 a_5840_15093.n2 a_5840_15093.t9 0.187648
R7964 a_5840_15093.n4 a_5840_15093.n3 0.0207092
R7965 a_5840_15093.n109 a_5840_15093.n4 0.0751921
R7966 a_5840_15093.n35 a_5840_15093.n34 0.0889741
R7967 a_5840_15093.n0 a_5840_15093.n4 0.318867
R7968 a_5840_15093.t9 a_5840_15093.n1 0.2981
R7969 a_5840_7613.t0 a_5840_7613.t1 25.621
R7970 a_22388_2038.t1 a_22388_2038.n1 21.2275
R7971 a_22388_2038.n1 a_22388_2038.t2 18.9805
R7972 a_22388_2038.n0 a_22388_2038.t5 17.5205
R7973 a_22388_2038.n0 a_22388_2038.t3 11.5588
R7974 a_22388_2038.n1 a_22388_2038.t4 11.4372
R7975 a_22388_2038.t1 a_22388_2038.t0 8.60523
R7976 a_22388_2038.t1 a_22388_2038.n0 8.27396
R7977 PLL_FREERUN.n75 PLL_FREERUN.t35 63.1691
R7978 PLL_FREERUN.t1 PLL_FREERUN.n26 58.6217
R7979 PLL_FREERUN.n9 PLL_FREERUN.t13 58.6217
R7980 PLL_FREERUN.n27 PLL_FREERUN.t1 55.3312
R7981 PLL_FREERUN.t13 PLL_FREERUN.n8 55.3312
R7982 PLL_FREERUN.n8 PLL_FREERUN.t14 39.8187
R7983 PLL_FREERUN.n9 PLL_FREERUN.t14 39.8187
R7984 PLL_FREERUN.n7 PLL_FREERUN.t32 39.8187
R7985 PLL_FREERUN.n10 PLL_FREERUN.t32 39.8187
R7986 PLL_FREERUN.n6 PLL_FREERUN.t5 39.8187
R7987 PLL_FREERUN.n11 PLL_FREERUN.t5 39.8187
R7988 PLL_FREERUN.n5 PLL_FREERUN.t24 39.8187
R7989 PLL_FREERUN.n12 PLL_FREERUN.t24 39.8187
R7990 PLL_FREERUN.n4 PLL_FREERUN.t9 39.8187
R7991 PLL_FREERUN.n13 PLL_FREERUN.t9 39.8187
R7992 PLL_FREERUN.n3 PLL_FREERUN.t27 39.8187
R7993 PLL_FREERUN.n14 PLL_FREERUN.t27 39.8187
R7994 PLL_FREERUN.n2 PLL_FREERUN.t15 39.8187
R7995 PLL_FREERUN.n15 PLL_FREERUN.t15 39.8187
R7996 PLL_FREERUN.n1 PLL_FREERUN.t3 39.8187
R7997 PLL_FREERUN.n16 PLL_FREERUN.t3 39.8187
R7998 PLL_FREERUN.t18 PLL_FREERUN.n0 39.8187
R7999 PLL_FREERUN.n17 PLL_FREERUN.t18 39.8187
R8000 PLL_FREERUN.n35 PLL_FREERUN.t37 39.8187
R8001 PLL_FREERUN.n18 PLL_FREERUN.t37 39.8187
R8002 PLL_FREERUN.n34 PLL_FREERUN.t23 39.8187
R8003 PLL_FREERUN.n19 PLL_FREERUN.t23 39.8187
R8004 PLL_FREERUN.n33 PLL_FREERUN.t40 39.8187
R8005 PLL_FREERUN.n20 PLL_FREERUN.t40 39.8187
R8006 PLL_FREERUN.n32 PLL_FREERUN.t30 39.8187
R8007 PLL_FREERUN.n21 PLL_FREERUN.t30 39.8187
R8008 PLL_FREERUN.n31 PLL_FREERUN.t4 39.8187
R8009 PLL_FREERUN.n22 PLL_FREERUN.t4 39.8187
R8010 PLL_FREERUN.n30 PLL_FREERUN.t34 39.8187
R8011 PLL_FREERUN.n23 PLL_FREERUN.t34 39.8187
R8012 PLL_FREERUN.n29 PLL_FREERUN.t7 39.8187
R8013 PLL_FREERUN.n24 PLL_FREERUN.t7 39.8187
R8014 PLL_FREERUN.n28 PLL_FREERUN.t25 39.8187
R8015 PLL_FREERUN.n25 PLL_FREERUN.t25 39.8187
R8016 PLL_FREERUN.n27 PLL_FREERUN.t11 39.8187
R8017 PLL_FREERUN.n26 PLL_FREERUN.t11 39.8187
R8018 PLL_FREERUN.n37 PLL_FREERUN.t38 37.0976
R8019 PLL_FREERUN.n47 PLL_FREERUN.t22 36.5005
R8020 PLL_FREERUN.t16 PLL_FREERUN.n64 36.5005
R8021 PLL_FREERUN.t22 PLL_FREERUN.n46 33.21
R8022 PLL_FREERUN.n65 PLL_FREERUN.t16 33.21
R8023 PLL_FREERUN.n48 PLL_FREERUN.n47 18.8035
R8024 PLL_FREERUN.n49 PLL_FREERUN.n48 18.8035
R8025 PLL_FREERUN.n50 PLL_FREERUN.n49 18.8035
R8026 PLL_FREERUN.n51 PLL_FREERUN.n50 18.8035
R8027 PLL_FREERUN.n52 PLL_FREERUN.n51 18.8035
R8028 PLL_FREERUN.n53 PLL_FREERUN.n52 18.8035
R8029 PLL_FREERUN.n54 PLL_FREERUN.n53 18.8035
R8030 PLL_FREERUN.n55 PLL_FREERUN.n54 18.8035
R8031 PLL_FREERUN.n56 PLL_FREERUN.n55 18.8035
R8032 PLL_FREERUN.n57 PLL_FREERUN.n56 18.8035
R8033 PLL_FREERUN.n58 PLL_FREERUN.n57 18.8035
R8034 PLL_FREERUN.n59 PLL_FREERUN.n58 18.8035
R8035 PLL_FREERUN.n60 PLL_FREERUN.n59 18.8035
R8036 PLL_FREERUN.n61 PLL_FREERUN.n60 18.8035
R8037 PLL_FREERUN.n62 PLL_FREERUN.n61 18.8035
R8038 PLL_FREERUN.n63 PLL_FREERUN.n62 18.8035
R8039 PLL_FREERUN.n64 PLL_FREERUN.n63 18.8035
R8040 PLL_FREERUN.n10 PLL_FREERUN.n9 18.8035
R8041 PLL_FREERUN.n11 PLL_FREERUN.n10 18.8035
R8042 PLL_FREERUN.n12 PLL_FREERUN.n11 18.8035
R8043 PLL_FREERUN.n13 PLL_FREERUN.n12 18.8035
R8044 PLL_FREERUN.n14 PLL_FREERUN.n13 18.8035
R8045 PLL_FREERUN.n15 PLL_FREERUN.n14 18.8035
R8046 PLL_FREERUN.n16 PLL_FREERUN.n15 18.8035
R8047 PLL_FREERUN.n17 PLL_FREERUN.n16 18.8035
R8048 PLL_FREERUN.n18 PLL_FREERUN.n17 18.8035
R8049 PLL_FREERUN.n19 PLL_FREERUN.n18 18.8035
R8050 PLL_FREERUN.n20 PLL_FREERUN.n19 18.8035
R8051 PLL_FREERUN.n21 PLL_FREERUN.n20 18.8035
R8052 PLL_FREERUN.n22 PLL_FREERUN.n21 18.8035
R8053 PLL_FREERUN.n23 PLL_FREERUN.n22 18.8035
R8054 PLL_FREERUN.n24 PLL_FREERUN.n23 18.8035
R8055 PLL_FREERUN.n25 PLL_FREERUN.n24 18.8035
R8056 PLL_FREERUN.n26 PLL_FREERUN.n25 18.8035
R8057 PLL_FREERUN.n65 PLL_FREERUN.t0 17.6975
R8058 PLL_FREERUN.n64 PLL_FREERUN.t0 17.6975
R8059 PLL_FREERUN.n66 PLL_FREERUN.t36 17.6975
R8060 PLL_FREERUN.n63 PLL_FREERUN.t36 17.6975
R8061 PLL_FREERUN.n67 PLL_FREERUN.t10 17.6975
R8062 PLL_FREERUN.n62 PLL_FREERUN.t10 17.6975
R8063 PLL_FREERUN.n68 PLL_FREERUN.t29 17.6975
R8064 PLL_FREERUN.n61 PLL_FREERUN.t29 17.6975
R8065 PLL_FREERUN.n69 PLL_FREERUN.t20 17.6975
R8066 PLL_FREERUN.n60 PLL_FREERUN.t20 17.6975
R8067 PLL_FREERUN.n70 PLL_FREERUN.t39 17.6975
R8068 PLL_FREERUN.n59 PLL_FREERUN.t39 17.6975
R8069 PLL_FREERUN.n71 PLL_FREERUN.t21 17.6975
R8070 PLL_FREERUN.n58 PLL_FREERUN.t21 17.6975
R8071 PLL_FREERUN.n72 PLL_FREERUN.t41 17.6975
R8072 PLL_FREERUN.n57 PLL_FREERUN.t41 17.6975
R8073 PLL_FREERUN.n73 PLL_FREERUN.t33 17.6975
R8074 PLL_FREERUN.n56 PLL_FREERUN.t33 17.6975
R8075 PLL_FREERUN.t8 PLL_FREERUN.n38 17.6975
R8076 PLL_FREERUN.n55 PLL_FREERUN.t8 17.6975
R8077 PLL_FREERUN.n39 PLL_FREERUN.t28 17.6975
R8078 PLL_FREERUN.n54 PLL_FREERUN.t28 17.6975
R8079 PLL_FREERUN.n40 PLL_FREERUN.t17 17.6975
R8080 PLL_FREERUN.n53 PLL_FREERUN.t17 17.6975
R8081 PLL_FREERUN.n41 PLL_FREERUN.t2 17.6975
R8082 PLL_FREERUN.n52 PLL_FREERUN.t2 17.6975
R8083 PLL_FREERUN.n42 PLL_FREERUN.t19 17.6975
R8084 PLL_FREERUN.n51 PLL_FREERUN.t19 17.6975
R8085 PLL_FREERUN.n43 PLL_FREERUN.t12 17.6975
R8086 PLL_FREERUN.n50 PLL_FREERUN.t12 17.6975
R8087 PLL_FREERUN.n44 PLL_FREERUN.t31 17.6975
R8088 PLL_FREERUN.n49 PLL_FREERUN.t31 17.6975
R8089 PLL_FREERUN.n45 PLL_FREERUN.t6 17.6975
R8090 PLL_FREERUN.n48 PLL_FREERUN.t6 17.6975
R8091 PLL_FREERUN.n46 PLL_FREERUN.t26 17.6975
R8092 PLL_FREERUN.n47 PLL_FREERUN.t26 17.6975
R8093 PLL_FREERUN.n46 PLL_FREERUN.n45 15.513
R8094 PLL_FREERUN.n45 PLL_FREERUN.n44 15.513
R8095 PLL_FREERUN.n44 PLL_FREERUN.n43 15.513
R8096 PLL_FREERUN.n43 PLL_FREERUN.n42 15.513
R8097 PLL_FREERUN.n42 PLL_FREERUN.n41 15.513
R8098 PLL_FREERUN.n41 PLL_FREERUN.n40 15.513
R8099 PLL_FREERUN.n40 PLL_FREERUN.n39 15.513
R8100 PLL_FREERUN.n39 PLL_FREERUN.n38 15.513
R8101 PLL_FREERUN.n73 PLL_FREERUN.n72 15.513
R8102 PLL_FREERUN.n72 PLL_FREERUN.n71 15.513
R8103 PLL_FREERUN.n71 PLL_FREERUN.n70 15.513
R8104 PLL_FREERUN.n70 PLL_FREERUN.n69 15.513
R8105 PLL_FREERUN.n69 PLL_FREERUN.n68 15.513
R8106 PLL_FREERUN.n68 PLL_FREERUN.n67 15.513
R8107 PLL_FREERUN.n67 PLL_FREERUN.n66 15.513
R8108 PLL_FREERUN.n66 PLL_FREERUN.n65 15.513
R8109 PLL_FREERUN.n8 PLL_FREERUN.n7 15.513
R8110 PLL_FREERUN.n7 PLL_FREERUN.n6 15.513
R8111 PLL_FREERUN.n6 PLL_FREERUN.n5 15.513
R8112 PLL_FREERUN.n5 PLL_FREERUN.n4 15.513
R8113 PLL_FREERUN.n4 PLL_FREERUN.n3 15.513
R8114 PLL_FREERUN.n3 PLL_FREERUN.n2 15.513
R8115 PLL_FREERUN.n2 PLL_FREERUN.n1 15.513
R8116 PLL_FREERUN.n1 PLL_FREERUN.n0 15.513
R8117 PLL_FREERUN.n35 PLL_FREERUN.n34 15.513
R8118 PLL_FREERUN.n34 PLL_FREERUN.n33 15.513
R8119 PLL_FREERUN.n33 PLL_FREERUN.n32 15.513
R8120 PLL_FREERUN.n32 PLL_FREERUN.n31 15.513
R8121 PLL_FREERUN.n31 PLL_FREERUN.n30 15.513
R8122 PLL_FREERUN.n30 PLL_FREERUN.n29 15.513
R8123 PLL_FREERUN.n29 PLL_FREERUN.n28 15.513
R8124 PLL_FREERUN.n28 PLL_FREERUN.n27 15.513
R8125 PLL_FREERUN.n74 PLL_FREERUN.n38 7.75675
R8126 PLL_FREERUN.n74 PLL_FREERUN.n73 7.75675
R8127 PLL_FREERUN.n36 PLL_FREERUN.n0 7.75675
R8128 PLL_FREERUN.n36 PLL_FREERUN.n35 7.75675
R8129 PLL_FREERUN.n37 PLL_FREERUN.n36 6.82995
R8130 PLL_FREERUN.n75 PLL_FREERUN.n74 6.82208
R8131 PLL_FREERUN PLL_FREERUN.n76 1.72963
R8132 PLL_FREERUN.n76 PLL_FREERUN.n75 0.77
R8133 PLL_FREERUN.n76 PLL_FREERUN.n37 0.487625
R8134 PLL_VCTRL.n29 PLL_VCTRL.n28 15.3005
R8135 PLL_VCTRL.n26 PLL_VCTRL.n25 15.3005
R8136 PLL_VCTRL.n23 PLL_VCTRL.n22 15.3005
R8137 PLL_VCTRL.n20 PLL_VCTRL.n19 15.3005
R8138 PLL_VCTRL.n17 PLL_VCTRL.n16 15.3005
R8139 PLL_VCTRL.n14 PLL_VCTRL.n13 15.3005
R8140 PLL_VCTRL.n11 PLL_VCTRL.n10 15.3005
R8141 PLL_VCTRL.n8 PLL_VCTRL.n7 15.3005
R8142 PLL_VCTRL.n5 PLL_VCTRL.n4 15.3005
R8143 PLL_VCTRL.n2 PLL_VCTRL.n1 15.3005
R8144 PLL_VCTRL.n29 PLL_VCTRL.n27 3.38042
R8145 PLL_VCTRL.n26 PLL_VCTRL.n24 3.38042
R8146 PLL_VCTRL.n23 PLL_VCTRL.n21 3.38042
R8147 PLL_VCTRL.n20 PLL_VCTRL.n18 3.38042
R8148 PLL_VCTRL.n17 PLL_VCTRL.n15 3.38042
R8149 PLL_VCTRL.n14 PLL_VCTRL.n12 3.38042
R8150 PLL_VCTRL.n11 PLL_VCTRL.n9 3.38042
R8151 PLL_VCTRL.n8 PLL_VCTRL.n6 3.38042
R8152 PLL_VCTRL.n5 PLL_VCTRL.n3 3.38042
R8153 PLL_VCTRL.n2 PLL_VCTRL.n0 3.38042
R8154 PLL_VCTRL PLL_VCTRL.n29 1.75994
R8155 PLL_VCTRL.n28 PLL_VCTRL.t15 1.6385
R8156 PLL_VCTRL.n28 PLL_VCTRL.t1 1.6385
R8157 PLL_VCTRL.n25 PLL_VCTRL.t17 1.6385
R8158 PLL_VCTRL.n25 PLL_VCTRL.t4 1.6385
R8159 PLL_VCTRL.n22 PLL_VCTRL.t12 1.6385
R8160 PLL_VCTRL.n22 PLL_VCTRL.t11 1.6385
R8161 PLL_VCTRL.n19 PLL_VCTRL.t3 1.6385
R8162 PLL_VCTRL.n19 PLL_VCTRL.t9 1.6385
R8163 PLL_VCTRL.n16 PLL_VCTRL.t5 1.6385
R8164 PLL_VCTRL.n16 PLL_VCTRL.t8 1.6385
R8165 PLL_VCTRL.n13 PLL_VCTRL.t18 1.6385
R8166 PLL_VCTRL.n13 PLL_VCTRL.t6 1.6385
R8167 PLL_VCTRL.n10 PLL_VCTRL.t14 1.6385
R8168 PLL_VCTRL.n10 PLL_VCTRL.t0 1.6385
R8169 PLL_VCTRL.n7 PLL_VCTRL.t16 1.6385
R8170 PLL_VCTRL.n7 PLL_VCTRL.t13 1.6385
R8171 PLL_VCTRL.n4 PLL_VCTRL.t7 1.6385
R8172 PLL_VCTRL.n4 PLL_VCTRL.t10 1.6385
R8173 PLL_VCTRL.n1 PLL_VCTRL.t2 1.6385
R8174 PLL_VCTRL.n1 PLL_VCTRL.t19 1.6385
R8175 PLL_VCTRL.n27 PLL_VCTRL.t25 0.607167
R8176 PLL_VCTRL.n27 PLL_VCTRL.t29 0.607167
R8177 PLL_VCTRL.n24 PLL_VCTRL.t38 0.607167
R8178 PLL_VCTRL.n24 PLL_VCTRL.t26 0.607167
R8179 PLL_VCTRL.n21 PLL_VCTRL.t27 0.607167
R8180 PLL_VCTRL.n21 PLL_VCTRL.t37 0.607167
R8181 PLL_VCTRL.n18 PLL_VCTRL.t30 0.607167
R8182 PLL_VCTRL.n18 PLL_VCTRL.t28 0.607167
R8183 PLL_VCTRL.n15 PLL_VCTRL.t24 0.607167
R8184 PLL_VCTRL.n15 PLL_VCTRL.t32 0.607167
R8185 PLL_VCTRL.n12 PLL_VCTRL.t35 0.607167
R8186 PLL_VCTRL.n12 PLL_VCTRL.t34 0.607167
R8187 PLL_VCTRL.n9 PLL_VCTRL.t20 0.607167
R8188 PLL_VCTRL.n9 PLL_VCTRL.t36 0.607167
R8189 PLL_VCTRL.n6 PLL_VCTRL.t23 0.607167
R8190 PLL_VCTRL.n6 PLL_VCTRL.t22 0.607167
R8191 PLL_VCTRL.n3 PLL_VCTRL.t33 0.607167
R8192 PLL_VCTRL.n3 PLL_VCTRL.t31 0.607167
R8193 PLL_VCTRL.n0 PLL_VCTRL.t21 0.607167
R8194 PLL_VCTRL.n0 PLL_VCTRL.t39 0.607167
R8195 PLL_VCTRL.n5 PLL_VCTRL.n2 0.0152683
R8196 PLL_VCTRL.n8 PLL_VCTRL.n5 0.0152683
R8197 PLL_VCTRL.n11 PLL_VCTRL.n8 0.0152683
R8198 PLL_VCTRL.n14 PLL_VCTRL.n11 0.0152683
R8199 PLL_VCTRL.n17 PLL_VCTRL.n14 0.0152683
R8200 PLL_VCTRL.n20 PLL_VCTRL.n17 0.0152683
R8201 PLL_VCTRL.n23 PLL_VCTRL.n20 0.0152683
R8202 PLL_VCTRL.n26 PLL_VCTRL.n23 0.0152683
R8203 PLL_VCTRL.n29 PLL_VCTRL.n26 0.0152683
R8204 DEBUG.n58 DEBUG.t80 29.6701
R8205 DEBUG.n28 DEBUG.t14 14.1508
R8206 DEBUG.n18 DEBUG.t19 14.1508
R8207 DEBUG.n57 DEBUG.t40 14.1508
R8208 DEBUG.n47 DEBUG.t66 14.1508
R8209 DEBUG.n27 DEBUG.n1 11.5047
R8210 DEBUG.n26 DEBUG.n3 11.5047
R8211 DEBUG.n25 DEBUG.n5 11.5047
R8212 DEBUG.n24 DEBUG.n7 11.5047
R8213 DEBUG.n23 DEBUG.n9 11.5047
R8214 DEBUG.n22 DEBUG.n11 11.5047
R8215 DEBUG.n21 DEBUG.n13 11.5047
R8216 DEBUG.n20 DEBUG.n15 11.5047
R8217 DEBUG.n19 DEBUG.n17 11.5047
R8218 DEBUG.n56 DEBUG.n30 11.5047
R8219 DEBUG.n55 DEBUG.n32 11.5047
R8220 DEBUG.n54 DEBUG.n34 11.5047
R8221 DEBUG.n53 DEBUG.n36 11.5047
R8222 DEBUG.n52 DEBUG.n38 11.5047
R8223 DEBUG.n51 DEBUG.n40 11.5047
R8224 DEBUG.n50 DEBUG.n42 11.5047
R8225 DEBUG.n49 DEBUG.n44 11.5047
R8226 DEBUG.n48 DEBUG.n46 11.5047
R8227 DEBUG.n28 DEBUG.t45 4.19837
R8228 DEBUG.n18 DEBUG.t59 4.19837
R8229 DEBUG.n57 DEBUG.t5 4.19837
R8230 DEBUG.n47 DEBUG.t29 4.19837
R8231 DEBUG.n27 DEBUG.n0 3.21837
R8232 DEBUG.n26 DEBUG.n2 3.21837
R8233 DEBUG.n25 DEBUG.n4 3.21837
R8234 DEBUG.n24 DEBUG.n6 3.21837
R8235 DEBUG.n23 DEBUG.n8 3.21837
R8236 DEBUG.n22 DEBUG.n10 3.21837
R8237 DEBUG.n21 DEBUG.n12 3.21837
R8238 DEBUG.n20 DEBUG.n14 3.21837
R8239 DEBUG.n19 DEBUG.n16 3.21837
R8240 DEBUG.n56 DEBUG.n29 3.21837
R8241 DEBUG.n55 DEBUG.n31 3.21837
R8242 DEBUG.n54 DEBUG.n33 3.21837
R8243 DEBUG.n53 DEBUG.n35 3.21837
R8244 DEBUG.n52 DEBUG.n37 3.21837
R8245 DEBUG.n51 DEBUG.n39 3.21837
R8246 DEBUG.n50 DEBUG.n41 3.21837
R8247 DEBUG.n49 DEBUG.n43 3.21837
R8248 DEBUG.n48 DEBUG.n45 3.21837
R8249 DEBUG.n58 DEBUG.n28 1.73975
R8250 DEBUG.n1 DEBUG.t13 1.6385
R8251 DEBUG.n1 DEBUG.t23 1.6385
R8252 DEBUG.n3 DEBUG.t10 1.6385
R8253 DEBUG.n3 DEBUG.t20 1.6385
R8254 DEBUG.n5 DEBUG.t17 1.6385
R8255 DEBUG.n5 DEBUG.t24 1.6385
R8256 DEBUG.n7 DEBUG.t18 1.6385
R8257 DEBUG.n7 DEBUG.t12 1.6385
R8258 DEBUG.n9 DEBUG.t22 1.6385
R8259 DEBUG.n9 DEBUG.t9 1.6385
R8260 DEBUG.n11 DEBUG.t6 1.6385
R8261 DEBUG.n11 DEBUG.t15 1.6385
R8262 DEBUG.n13 DEBUG.t7 1.6385
R8263 DEBUG.n13 DEBUG.t16 1.6385
R8264 DEBUG.n15 DEBUG.t11 1.6385
R8265 DEBUG.n15 DEBUG.t21 1.6385
R8266 DEBUG.n17 DEBUG.t8 1.6385
R8267 DEBUG.n17 DEBUG.t25 1.6385
R8268 DEBUG.n30 DEBUG.t41 1.6385
R8269 DEBUG.n30 DEBUG.t49 1.6385
R8270 DEBUG.n32 DEBUG.t72 1.6385
R8271 DEBUG.n32 DEBUG.t79 1.6385
R8272 DEBUG.n34 DEBUG.t43 1.6385
R8273 DEBUG.n34 DEBUG.t58 1.6385
R8274 DEBUG.n36 DEBUG.t46 1.6385
R8275 DEBUG.n36 DEBUG.t67 1.6385
R8276 DEBUG.n38 DEBUG.t62 1.6385
R8277 DEBUG.n38 DEBUG.t51 1.6385
R8278 DEBUG.n40 DEBUG.t70 1.6385
R8279 DEBUG.n40 DEBUG.t65 1.6385
R8280 DEBUG.n42 DEBUG.t60 1.6385
R8281 DEBUG.n42 DEBUG.t71 1.6385
R8282 DEBUG.n44 DEBUG.t50 1.6385
R8283 DEBUG.n44 DEBUG.t73 1.6385
R8284 DEBUG.n46 DEBUG.t56 1.6385
R8285 DEBUG.n46 DEBUG.t44 1.6385
R8286 DEBUG.n0 DEBUG.t78 0.607167
R8287 DEBUG.n0 DEBUG.t68 0.607167
R8288 DEBUG.n2 DEBUG.t63 0.607167
R8289 DEBUG.n2 DEBUG.t48 0.607167
R8290 DEBUG.n4 DEBUG.t47 0.607167
R8291 DEBUG.n4 DEBUG.t42 0.607167
R8292 DEBUG.n6 DEBUG.t75 0.607167
R8293 DEBUG.n6 DEBUG.t74 0.607167
R8294 DEBUG.n8 DEBUG.t69 0.607167
R8295 DEBUG.n8 DEBUG.t52 0.607167
R8296 DEBUG.n10 DEBUG.t64 0.607167
R8297 DEBUG.n10 DEBUG.t61 0.607167
R8298 DEBUG.n12 DEBUG.t57 0.607167
R8299 DEBUG.n12 DEBUG.t55 0.607167
R8300 DEBUG.n14 DEBUG.t76 0.607167
R8301 DEBUG.n14 DEBUG.t77 0.607167
R8302 DEBUG.n16 DEBUG.t54 0.607167
R8303 DEBUG.n16 DEBUG.t53 0.607167
R8304 DEBUG.n29 DEBUG.t4 0.607167
R8305 DEBUG.n29 DEBUG.t33 0.607167
R8306 DEBUG.n31 DEBUG.t26 0.607167
R8307 DEBUG.n31 DEBUG.t0 0.607167
R8308 DEBUG.n33 DEBUG.t38 0.607167
R8309 DEBUG.n33 DEBUG.t35 0.607167
R8310 DEBUG.n35 DEBUG.t3 0.607167
R8311 DEBUG.n35 DEBUG.t28 0.607167
R8312 DEBUG.n37 DEBUG.t2 0.607167
R8313 DEBUG.n37 DEBUG.t31 0.607167
R8314 DEBUG.n39 DEBUG.t1 0.607167
R8315 DEBUG.n39 DEBUG.t30 0.607167
R8316 DEBUG.n41 DEBUG.t34 0.607167
R8317 DEBUG.n41 DEBUG.t27 0.607167
R8318 DEBUG.n43 DEBUG.t32 0.607167
R8319 DEBUG.n43 DEBUG.t39 0.607167
R8320 DEBUG.n45 DEBUG.t36 0.607167
R8321 DEBUG.n45 DEBUG.t37 0.607167
R8322 DEBUG.n58 DEBUG.n57 0.21245
R8323 DEBUG.n28 DEBUG.n27 0.1679
R8324 DEBUG.n19 DEBUG.n18 0.1679
R8325 DEBUG.n57 DEBUG.n56 0.1679
R8326 DEBUG.n48 DEBUG.n47 0.1679
R8327 DEBUG.n27 DEBUG.n26 0.1535
R8328 DEBUG.n26 DEBUG.n25 0.1535
R8329 DEBUG.n25 DEBUG.n24 0.1535
R8330 DEBUG.n24 DEBUG.n23 0.1535
R8331 DEBUG.n23 DEBUG.n22 0.1535
R8332 DEBUG.n22 DEBUG.n21 0.1535
R8333 DEBUG.n21 DEBUG.n20 0.1535
R8334 DEBUG.n20 DEBUG.n19 0.1535
R8335 DEBUG.n56 DEBUG.n55 0.1535
R8336 DEBUG.n55 DEBUG.n54 0.1535
R8337 DEBUG.n54 DEBUG.n53 0.1535
R8338 DEBUG.n53 DEBUG.n52 0.1535
R8339 DEBUG.n52 DEBUG.n51 0.1535
R8340 DEBUG.n51 DEBUG.n50 0.1535
R8341 DEBUG.n50 DEBUG.n49 0.1535
R8342 DEBUG.n49 DEBUG.n48 0.1535
R8343 DEBUG DEBUG.n58 0.02255
R8344 PLL_DISABLE.n9 PLL_DISABLE.t7 58.6217
R8345 PLL_DISABLE.t19 PLL_DISABLE.n26 58.6217
R8346 PLL_DISABLE.t7 PLL_DISABLE.n8 55.3312
R8347 PLL_DISABLE.n27 PLL_DISABLE.t19 55.3312
R8348 PLL_DISABLE.n27 PLL_DISABLE.t1 39.8187
R8349 PLL_DISABLE.n26 PLL_DISABLE.t1 39.8187
R8350 PLL_DISABLE.n28 PLL_DISABLE.t17 39.8187
R8351 PLL_DISABLE.n25 PLL_DISABLE.t17 39.8187
R8352 PLL_DISABLE.n29 PLL_DISABLE.t4 39.8187
R8353 PLL_DISABLE.n24 PLL_DISABLE.t4 39.8187
R8354 PLL_DISABLE.n30 PLL_DISABLE.t11 39.8187
R8355 PLL_DISABLE.n23 PLL_DISABLE.t11 39.8187
R8356 PLL_DISABLE.n31 PLL_DISABLE.t34 39.8187
R8357 PLL_DISABLE.n22 PLL_DISABLE.t34 39.8187
R8358 PLL_DISABLE.n32 PLL_DISABLE.t14 39.8187
R8359 PLL_DISABLE.n21 PLL_DISABLE.t14 39.8187
R8360 PLL_DISABLE.n33 PLL_DISABLE.t15 39.8187
R8361 PLL_DISABLE.n20 PLL_DISABLE.t15 39.8187
R8362 PLL_DISABLE.n34 PLL_DISABLE.t2 39.8187
R8363 PLL_DISABLE.n19 PLL_DISABLE.t2 39.8187
R8364 PLL_DISABLE.n35 PLL_DISABLE.t21 39.8187
R8365 PLL_DISABLE.n18 PLL_DISABLE.t21 39.8187
R8366 PLL_DISABLE.t30 PLL_DISABLE.n0 39.8187
R8367 PLL_DISABLE.n17 PLL_DISABLE.t30 39.8187
R8368 PLL_DISABLE.n1 PLL_DISABLE.t12 39.8187
R8369 PLL_DISABLE.n16 PLL_DISABLE.t12 39.8187
R8370 PLL_DISABLE.n2 PLL_DISABLE.t36 39.8187
R8371 PLL_DISABLE.n15 PLL_DISABLE.t36 39.8187
R8372 PLL_DISABLE.n3 PLL_DISABLE.t26 39.8187
R8373 PLL_DISABLE.n14 PLL_DISABLE.t26 39.8187
R8374 PLL_DISABLE.n4 PLL_DISABLE.t0 39.8187
R8375 PLL_DISABLE.n13 PLL_DISABLE.t0 39.8187
R8376 PLL_DISABLE.n5 PLL_DISABLE.t16 39.8187
R8377 PLL_DISABLE.n12 PLL_DISABLE.t16 39.8187
R8378 PLL_DISABLE.n6 PLL_DISABLE.t3 39.8187
R8379 PLL_DISABLE.n11 PLL_DISABLE.t3 39.8187
R8380 PLL_DISABLE.n7 PLL_DISABLE.t9 39.8187
R8381 PLL_DISABLE.n10 PLL_DISABLE.t9 39.8187
R8382 PLL_DISABLE.n8 PLL_DISABLE.t31 39.8187
R8383 PLL_DISABLE.n9 PLL_DISABLE.t31 39.8187
R8384 PLL_DISABLE.n10 PLL_DISABLE.n9 18.8035
R8385 PLL_DISABLE.n11 PLL_DISABLE.n10 18.8035
R8386 PLL_DISABLE.n12 PLL_DISABLE.n11 18.8035
R8387 PLL_DISABLE.n13 PLL_DISABLE.n12 18.8035
R8388 PLL_DISABLE.n14 PLL_DISABLE.n13 18.8035
R8389 PLL_DISABLE.n15 PLL_DISABLE.n14 18.8035
R8390 PLL_DISABLE.n16 PLL_DISABLE.n15 18.8035
R8391 PLL_DISABLE.n17 PLL_DISABLE.n16 18.8035
R8392 PLL_DISABLE.n18 PLL_DISABLE.n17 18.8035
R8393 PLL_DISABLE.n19 PLL_DISABLE.n18 18.8035
R8394 PLL_DISABLE.n20 PLL_DISABLE.n19 18.8035
R8395 PLL_DISABLE.n21 PLL_DISABLE.n20 18.8035
R8396 PLL_DISABLE.n22 PLL_DISABLE.n21 18.8035
R8397 PLL_DISABLE.n23 PLL_DISABLE.n22 18.8035
R8398 PLL_DISABLE.n24 PLL_DISABLE.n23 18.8035
R8399 PLL_DISABLE.n25 PLL_DISABLE.n24 18.8035
R8400 PLL_DISABLE.n26 PLL_DISABLE.n25 18.8035
R8401 PLL_DISABLE.n8 PLL_DISABLE.n7 15.513
R8402 PLL_DISABLE.n7 PLL_DISABLE.n6 15.513
R8403 PLL_DISABLE.n6 PLL_DISABLE.n5 15.513
R8404 PLL_DISABLE.n5 PLL_DISABLE.n4 15.513
R8405 PLL_DISABLE.n4 PLL_DISABLE.n3 15.513
R8406 PLL_DISABLE.n3 PLL_DISABLE.n2 15.513
R8407 PLL_DISABLE.n2 PLL_DISABLE.n1 15.513
R8408 PLL_DISABLE.n1 PLL_DISABLE.n0 15.513
R8409 PLL_DISABLE.n35 PLL_DISABLE.n34 15.513
R8410 PLL_DISABLE.n34 PLL_DISABLE.n33 15.513
R8411 PLL_DISABLE.n33 PLL_DISABLE.n32 15.513
R8412 PLL_DISABLE.n32 PLL_DISABLE.n31 15.513
R8413 PLL_DISABLE.n31 PLL_DISABLE.n30 15.513
R8414 PLL_DISABLE.n30 PLL_DISABLE.n29 15.513
R8415 PLL_DISABLE.n29 PLL_DISABLE.n28 15.513
R8416 PLL_DISABLE.n28 PLL_DISABLE.n27 15.513
R8417 PLL_DISABLE.n42 PLL_DISABLE.t13 15.4765
R8418 PLL_DISABLE.n43 PLL_DISABLE.t25 15.4765
R8419 PLL_DISABLE.n45 PLL_DISABLE.t6 15.4765
R8420 PLL_DISABLE.n46 PLL_DISABLE.t28 15.4765
R8421 PLL_DISABLE.n47 PLL_DISABLE.t8 15.4765
R8422 PLL_DISABLE.n48 PLL_DISABLE.t18 15.4765
R8423 PLL_DISABLE.n40 PLL_DISABLE.t20 15.4765
R8424 PLL_DISABLE.n41 PLL_DISABLE.t10 15.4765
R8425 PLL_DISABLE.n42 PLL_DISABLE.t33 13.7488
R8426 PLL_DISABLE.n43 PLL_DISABLE.t32 13.7488
R8427 PLL_DISABLE.n45 PLL_DISABLE.t24 13.7488
R8428 PLL_DISABLE.n46 PLL_DISABLE.t35 13.7488
R8429 PLL_DISABLE.n47 PLL_DISABLE.t27 13.7488
R8430 PLL_DISABLE.n48 PLL_DISABLE.t22 13.7488
R8431 PLL_DISABLE.n40 PLL_DISABLE.t23 13.7488
R8432 PLL_DISABLE.n41 PLL_DISABLE.t29 13.7488
R8433 PLL_DISABLE.n43 PLL_DISABLE.n42 10.5449
R8434 PLL_DISABLE.n46 PLL_DISABLE.n45 10.5449
R8435 PLL_DISABLE.n47 PLL_DISABLE.n46 10.5449
R8436 PLL_DISABLE.n48 PLL_DISABLE.n47 10.5449
R8437 PLL_DISABLE.n41 PLL_DISABLE.n40 10.5449
R8438 PLL_DISABLE.n38 PLL_DISABLE.n37 9.0005
R8439 PLL_DISABLE.n45 PLL_DISABLE.n44 8.41578
R8440 PLL_DISABLE.n38 PLL_DISABLE.n36 7.89365
R8441 PLL_DISABLE.n36 PLL_DISABLE.n0 7.75675
R8442 PLL_DISABLE.n36 PLL_DISABLE.n35 7.75675
R8443 PLL_DISABLE.n37 PLL_DISABLE.t37 6.54431
R8444 PLL_DISABLE.n49 PLL_DISABLE.n48 6.388
R8445 PLL_DISABLE.n50 PLL_DISABLE.n49 6.00626
R8446 PLL_DISABLE.n44 PLL_DISABLE.n39 5.9799
R8447 PLL_DISABLE.n37 PLL_DISABLE.t5 5.35834
R8448 PLL_DISABLE PLL_DISABLE.n50 4.98875
R8449 PLL_DISABLE.n49 PLL_DISABLE.n41 4.15744
R8450 PLL_DISABLE.n44 PLL_DISABLE.n43 2.12967
R8451 PLL_DISABLE.n50 PLL_DISABLE.n39 1.96025
R8452 PLL_DISABLE.n39 PLL_DISABLE.n38 0.4235
R8453 a_n15085_2072.n30 a_n15085_2072.n36 17.042
R8454 a_n15085_2072.n1 a_n15085_2072.n49 17.042
R8455 a_n15085_2072.n32 a_n15085_2072.n48 17.042
R8456 a_n15085_2072.n23 a_n15085_2072.n47 17.042
R8457 a_n15085_2072.n27 a_n15085_2072.n45 17.042
R8458 a_n15085_2072.n26 a_n15085_2072.n44 17.042
R8459 a_n15085_2072.n34 a_n15085_2072.n42 17.042
R8460 a_n15085_2072.n31 a_n15085_2072.n40 17.042
R8461 a_n15085_2072.n4 a_n15085_2072.n39 17.042
R8462 a_n15085_2072.n29 a_n15085_2072.n37 17.042
R8463 a_n15085_2072.n6 a_n15085_2072.t20 14.8576
R8464 a_n15085_2072.n25 a_n15085_2072.n12 0.74518
R8465 a_n15085_2072.n13 a_n15085_2072.n12 1.12134
R8466 a_n15085_2072.n14 a_n15085_2072.n12 0.637352
R8467 a_n15085_2072.n15 a_n15085_2072.n12 0.744654
R8468 a_n15085_2072.n16 a_n15085_2072.n12 0.744654
R8469 a_n15085_2072.n17 a_n15085_2072.n12 0.744654
R8470 a_n15085_2072.n18 a_n15085_2072.n12 0.744654
R8471 a_n15085_2072.n19 a_n15085_2072.n12 0.744654
R8472 a_n15085_2072.n20 a_n15085_2072.n12 0.744654
R8473 a_n15085_2072.n8 a_n15085_2072.n12 0.744654
R8474 a_n15085_2072.n11 a_n15085_2072.n12 0.397292
R8475 a_n15085_2072.n1 a_n15085_2072.n50 3.38042
R8476 a_n15085_2072.n32 a_n15085_2072.n51 3.38042
R8477 a_n15085_2072.n23 a_n15085_2072.n53 3.38042
R8478 a_n15085_2072.n27 a_n15085_2072.n46 3.38042
R8479 a_n15085_2072.n26 a_n15085_2072.n59 3.38042
R8480 a_n15085_2072.n34 a_n15085_2072.n43 3.38042
R8481 a_n15085_2072.n31 a_n15085_2072.n41 3.38042
R8482 a_n15085_2072.n4 a_n15085_2072.n65 3.38042
R8483 a_n15085_2072.n29 a_n15085_2072.n38 3.38042
R8484 a_n15085_2072.n67 a_n15085_2072.n30 3.38042
R8485 a_n15085_2072.n66 a_n15085_2072.n25 0.0136025
R8486 a_n15085_2072.n12 a_n15085_2072.n7 0.893651
R8487 a_n15085_2072.n11 a_n15085_2072.n0 0.773659
R8488 a_n15085_2072.n36 a_n15085_2072.t24 1.6385
R8489 a_n15085_2072.n36 a_n15085_2072.t34 1.6385
R8490 a_n15085_2072.n49 a_n15085_2072.t39 1.6385
R8491 a_n15085_2072.n49 a_n15085_2072.t29 1.6385
R8492 a_n15085_2072.n48 a_n15085_2072.t37 1.6385
R8493 a_n15085_2072.n48 a_n15085_2072.t27 1.6385
R8494 a_n15085_2072.n47 a_n15085_2072.t33 1.6385
R8495 a_n15085_2072.n47 a_n15085_2072.t31 1.6385
R8496 a_n15085_2072.n45 a_n15085_2072.t28 1.6385
R8497 a_n15085_2072.n45 a_n15085_2072.t36 1.6385
R8498 a_n15085_2072.n44 a_n15085_2072.t35 1.6385
R8499 a_n15085_2072.n44 a_n15085_2072.t32 1.6385
R8500 a_n15085_2072.n42 a_n15085_2072.t30 1.6385
R8501 a_n15085_2072.n42 a_n15085_2072.t25 1.6385
R8502 a_n15085_2072.n40 a_n15085_2072.t40 1.6385
R8503 a_n15085_2072.n40 a_n15085_2072.t23 1.6385
R8504 a_n15085_2072.n39 a_n15085_2072.t26 1.6385
R8505 a_n15085_2072.n39 a_n15085_2072.t38 1.6385
R8506 a_n15085_2072.n37 a_n15085_2072.t21 1.6385
R8507 a_n15085_2072.n37 a_n15085_2072.t22 1.6385
R8508 a_n15085_2072.n28 a_n15085_2072.n66 1.5005
R8509 a_n15085_2072.n13 a_n15085_2072.n5 0.0133805
R8510 a_n15085_2072.n4 a_n15085_2072.n5 0.74481
R8511 a_n15085_2072.n14 a_n15085_2072.n3 1.5005
R8512 a_n15085_2072.n31 a_n15085_2072.n64 1.5005
R8513 a_n15085_2072.n15 a_n15085_2072.n63 1.5005
R8514 a_n15085_2072.n62 a_n15085_2072.n61 1.5005
R8515 a_n15085_2072.n16 a_n15085_2072.n34 1.5005
R8516 a_n15085_2072.n33 a_n15085_2072.n60 1.5005
R8517 a_n15085_2072.n17 a_n15085_2072.n21 1.5005
R8518 a_n15085_2072.n26 a_n15085_2072.n58 1.5005
R8519 a_n15085_2072.n18 a_n15085_2072.n22 1.5005
R8520 a_n15085_2072.n27 a_n15085_2072.n57 1.5005
R8521 a_n15085_2072.n19 a_n15085_2072.n56 1.5005
R8522 a_n15085_2072.n55 a_n15085_2072.n54 1.5005
R8523 a_n15085_2072.n20 a_n15085_2072.n23 1.5005
R8524 a_n15085_2072.n35 a_n15085_2072.n52 1.5005
R8525 a_n15085_2072.n8 a_n15085_2072.n24 1.5005
R8526 a_n15085_2072.n32 a_n15085_2072.n10 0.012441
R8527 a_n15085_2072.n9 a_n15085_2072.n10 0.745279
R8528 a_n15085_2072.n2 a_n15085_2072.n7 0.0133857
R8529 a_n15085_2072.n2 a_n15085_2072.n1 0.744807
R8530 a_n15085_2072.n50 a_n15085_2072.t15 0.607167
R8531 a_n15085_2072.n50 a_n15085_2072.t6 0.607167
R8532 a_n15085_2072.n51 a_n15085_2072.t17 0.607167
R8533 a_n15085_2072.n51 a_n15085_2072.t2 0.607167
R8534 a_n15085_2072.n53 a_n15085_2072.t0 0.607167
R8535 a_n15085_2072.n53 a_n15085_2072.t4 0.607167
R8536 a_n15085_2072.n46 a_n15085_2072.t1 0.607167
R8537 a_n15085_2072.n46 a_n15085_2072.t8 0.607167
R8538 a_n15085_2072.n59 a_n15085_2072.t18 0.607167
R8539 a_n15085_2072.n59 a_n15085_2072.t9 0.607167
R8540 a_n15085_2072.n43 a_n15085_2072.t5 0.607167
R8541 a_n15085_2072.n43 a_n15085_2072.t10 0.607167
R8542 a_n15085_2072.n41 a_n15085_2072.t7 0.607167
R8543 a_n15085_2072.n41 a_n15085_2072.t14 0.607167
R8544 a_n15085_2072.n65 a_n15085_2072.t3 0.607167
R8545 a_n15085_2072.n65 a_n15085_2072.t16 0.607167
R8546 a_n15085_2072.n38 a_n15085_2072.t12 0.607167
R8547 a_n15085_2072.n38 a_n15085_2072.t11 0.607167
R8548 a_n15085_2072.n67 a_n15085_2072.t13 0.607167
R8549 a_n15085_2072.t19 a_n15085_2072.n67 0.607167
R8550 a_n15085_2072.n12 a_n15085_2072.n6 0.128009
R8551 a_n15085_2072.n6 a_n15085_2072.t47 0.063
R8552 a_n15085_2072.n6 a_n15085_2072.t50 0.063
R8553 a_n15085_2072.n6 a_n15085_2072.t49 0.063
R8554 a_n15085_2072.n6 a_n15085_2072.t44 0.063
R8555 a_n15085_2072.n6 a_n15085_2072.t41 0.063
R8556 a_n15085_2072.n6 a_n15085_2072.t45 0.063
R8557 a_n15085_2072.n6 a_n15085_2072.t48 0.063
R8558 a_n15085_2072.n6 a_n15085_2072.t43 0.063
R8559 a_n15085_2072.n6 a_n15085_2072.t42 0.063
R8560 a_n15085_2072.n30 a_n15085_2072.n0 0.01631
R8561 a_n15085_2072.n29 a_n15085_2072.n28 0.0313678
R8562 a_n15085_2072.n66 a_n15085_2072.n13 0.0235579
R8563 a_n15085_2072.n4 a_n15085_2072.n3 0.0235579
R8564 a_n15085_2072.n3 a_n15085_2072.n31 0.0235579
R8565 a_n15085_2072.n63 a_n15085_2072.n62 0.0235579
R8566 a_n15085_2072.n34 a_n15085_2072.n33 0.0235579
R8567 a_n15085_2072.n33 a_n15085_2072.n21 0.0235579
R8568 a_n15085_2072.n26 a_n15085_2072.n22 0.0235579
R8569 a_n15085_2072.n22 a_n15085_2072.n27 0.0235579
R8570 a_n15085_2072.n56 a_n15085_2072.n55 0.0235579
R8571 a_n15085_2072.n55 a_n15085_2072.n23 0.0235579
R8572 a_n15085_2072.n35 a_n15085_2072.n24 0.0235579
R8573 a_n15085_2072.n1 a_n15085_2072.n0 0.0393019
R8574 a_n15085_2072.n23 a_n15085_2072.n35 0.0235579
R8575 a_n15085_2072.n62 a_n15085_2072.n34 0.0235579
R8576 a_n15085_2072.n24 a_n15085_2072.n32 0.0235579
R8577 a_n15085_2072.n63 a_n15085_2072.n31 0.0235579
R8578 a_n15085_2072.n56 a_n15085_2072.n27 0.0235579
R8579 a_n15085_2072.n21 a_n15085_2072.n26 0.0235579
R8580 a_n15085_2072.n25 a_n15085_2072.n29 1.51326
R8581 a_n15085_2072.n6 a_n15085_2072.t46 0.0839524
R8582 a_n15085_2072.n10 a_n15085_2072.n1 0.0585567
R8583 a_n15085_2072.n28 a_n15085_2072.n4 0.0466157
R8584 a_n15085_2072.n9 a_n15085_2072.n8 0.0428732
R8585 a_n15085_2072.n9 a_n15085_2072.n7 0.0338789
R8586 a_n15085_2072.n52 a_n15085_2072.n20 0.0263872
R8587 a_n15085_2072.n54 a_n15085_2072.n19 0.0263872
R8588 a_n15085_2072.n57 a_n15085_2072.n18 0.0263872
R8589 a_n15085_2072.n58 a_n15085_2072.n17 0.0263872
R8590 a_n15085_2072.n60 a_n15085_2072.n16 0.0263872
R8591 a_n15085_2072.n61 a_n15085_2072.n15 0.0263872
R8592 a_n15085_2072.n64 a_n15085_2072.n14 0.0263744
R8593 a_n15085_2072.n2 a_n15085_2072.n11 0.0299138
R8594 a_n15085_2072.n52 a_n15085_2072.n8 0.0254776
R8595 a_n15085_2072.n54 a_n15085_2072.n20 0.0254776
R8596 a_n15085_2072.n57 a_n15085_2072.n19 0.0254776
R8597 a_n15085_2072.n58 a_n15085_2072.n18 0.0254776
R8598 a_n15085_2072.n60 a_n15085_2072.n17 0.0254776
R8599 a_n15085_2072.n61 a_n15085_2072.n16 0.0254776
R8600 a_n15085_2072.n64 a_n15085_2072.n15 0.0254776
R8601 a_n15085_2072.n14 a_n15085_2072.n5 0.0393129
R8602 a_n558_2704.n3 a_n558_2704.t8 39.434
R8603 a_n558_2704.n0 a_n558_2704.t6 39.3425
R8604 a_n558_2704.n0 a_n558_2704.t7 29.4555
R8605 a_n558_2704.n3 a_n558_2704.t5 29.3205
R8606 a_n558_2704.n1 a_n558_2704.t4 28.7301
R8607 a_n558_2704.n1 a_n558_2704.t3 18.7615
R8608 a_n558_2704.n2 a_n558_2704.t1 13.7342
R8609 a_n558_2704.n1 a_n558_2704.t2 13.5055
R8610 a_n558_2704.n0 a_n558_2704.n1 9.0247
R8611 a_n558_2704.n2 a_n558_2704.n3 7.96025
R8612 a_n558_2704.t0 a_n558_2704.n2 6.3271
R8613 a_n558_2704.n2 a_n558_2704.n0 1.39825
R8614 a_n17351_68.t21 a_n17351_68.n64 58.6217
R8615 a_n17351_68.n47 a_n17351_68.t34 58.6217
R8616 a_n17351_68.n65 a_n17351_68.t21 55.3312
R8617 a_n17351_68.t34 a_n17351_68.n46 55.3312
R8618 a_n17351_68.n46 a_n17351_68.t12 39.8187
R8619 a_n17351_68.n47 a_n17351_68.t12 39.8187
R8620 a_n17351_68.n45 a_n17351_68.t8 39.8187
R8621 a_n17351_68.n48 a_n17351_68.t8 39.8187
R8622 a_n17351_68.n44 a_n17351_68.t3 39.8187
R8623 a_n17351_68.n49 a_n17351_68.t3 39.8187
R8624 a_n17351_68.n43 a_n17351_68.t40 39.8187
R8625 a_n17351_68.n50 a_n17351_68.t40 39.8187
R8626 a_n17351_68.n42 a_n17351_68.t39 39.8187
R8627 a_n17351_68.n51 a_n17351_68.t39 39.8187
R8628 a_n17351_68.n41 a_n17351_68.t37 39.8187
R8629 a_n17351_68.n52 a_n17351_68.t37 39.8187
R8630 a_n17351_68.n40 a_n17351_68.t15 39.8187
R8631 a_n17351_68.n53 a_n17351_68.t15 39.8187
R8632 a_n17351_68.n39 a_n17351_68.t14 39.8187
R8633 a_n17351_68.n54 a_n17351_68.t14 39.8187
R8634 a_n17351_68.t9 a_n17351_68.n38 39.8187
R8635 a_n17351_68.n55 a_n17351_68.t9 39.8187
R8636 a_n17351_68.n73 a_n17351_68.t5 39.8187
R8637 a_n17351_68.n56 a_n17351_68.t5 39.8187
R8638 a_n17351_68.n72 a_n17351_68.t4 39.8187
R8639 a_n17351_68.n57 a_n17351_68.t4 39.8187
R8640 a_n17351_68.n71 a_n17351_68.t41 39.8187
R8641 a_n17351_68.n58 a_n17351_68.t41 39.8187
R8642 a_n17351_68.n70 a_n17351_68.t19 39.8187
R8643 a_n17351_68.n59 a_n17351_68.t19 39.8187
R8644 a_n17351_68.n69 a_n17351_68.t17 39.8187
R8645 a_n17351_68.n60 a_n17351_68.t17 39.8187
R8646 a_n17351_68.n68 a_n17351_68.t16 39.8187
R8647 a_n17351_68.n61 a_n17351_68.t16 39.8187
R8648 a_n17351_68.n67 a_n17351_68.t11 39.8187
R8649 a_n17351_68.n62 a_n17351_68.t11 39.8187
R8650 a_n17351_68.n66 a_n17351_68.t7 39.8187
R8651 a_n17351_68.n63 a_n17351_68.t7 39.8187
R8652 a_n17351_68.n65 a_n17351_68.t6 39.8187
R8653 a_n17351_68.n64 a_n17351_68.t6 39.8187
R8654 a_n17351_68.n10 a_n17351_68.t35 36.5005
R8655 a_n17351_68.t27 a_n17351_68.n27 36.5005
R8656 a_n17351_68.t35 a_n17351_68.n9 33.21
R8657 a_n17351_68.n28 a_n17351_68.t27 33.21
R8658 a_n17351_68.n11 a_n17351_68.n10 18.8035
R8659 a_n17351_68.n12 a_n17351_68.n11 18.8035
R8660 a_n17351_68.n13 a_n17351_68.n12 18.8035
R8661 a_n17351_68.n14 a_n17351_68.n13 18.8035
R8662 a_n17351_68.n15 a_n17351_68.n14 18.8035
R8663 a_n17351_68.n16 a_n17351_68.n15 18.8035
R8664 a_n17351_68.n17 a_n17351_68.n16 18.8035
R8665 a_n17351_68.n18 a_n17351_68.n17 18.8035
R8666 a_n17351_68.n19 a_n17351_68.n18 18.8035
R8667 a_n17351_68.n20 a_n17351_68.n19 18.8035
R8668 a_n17351_68.n21 a_n17351_68.n20 18.8035
R8669 a_n17351_68.n22 a_n17351_68.n21 18.8035
R8670 a_n17351_68.n23 a_n17351_68.n22 18.8035
R8671 a_n17351_68.n24 a_n17351_68.n23 18.8035
R8672 a_n17351_68.n25 a_n17351_68.n24 18.8035
R8673 a_n17351_68.n26 a_n17351_68.n25 18.8035
R8674 a_n17351_68.n27 a_n17351_68.n26 18.8035
R8675 a_n17351_68.n48 a_n17351_68.n47 18.8035
R8676 a_n17351_68.n49 a_n17351_68.n48 18.8035
R8677 a_n17351_68.n50 a_n17351_68.n49 18.8035
R8678 a_n17351_68.n51 a_n17351_68.n50 18.8035
R8679 a_n17351_68.n52 a_n17351_68.n51 18.8035
R8680 a_n17351_68.n53 a_n17351_68.n52 18.8035
R8681 a_n17351_68.n54 a_n17351_68.n53 18.8035
R8682 a_n17351_68.n55 a_n17351_68.n54 18.8035
R8683 a_n17351_68.n56 a_n17351_68.n55 18.8035
R8684 a_n17351_68.n57 a_n17351_68.n56 18.8035
R8685 a_n17351_68.n58 a_n17351_68.n57 18.8035
R8686 a_n17351_68.n59 a_n17351_68.n58 18.8035
R8687 a_n17351_68.n60 a_n17351_68.n59 18.8035
R8688 a_n17351_68.n61 a_n17351_68.n60 18.8035
R8689 a_n17351_68.n62 a_n17351_68.n61 18.8035
R8690 a_n17351_68.n63 a_n17351_68.n62 18.8035
R8691 a_n17351_68.n64 a_n17351_68.n63 18.8035
R8692 a_n17351_68.n28 a_n17351_68.t33 17.6975
R8693 a_n17351_68.n27 a_n17351_68.t33 17.6975
R8694 a_n17351_68.n29 a_n17351_68.t18 17.6975
R8695 a_n17351_68.n26 a_n17351_68.t18 17.6975
R8696 a_n17351_68.n30 a_n17351_68.t31 17.6975
R8697 a_n17351_68.n25 a_n17351_68.t31 17.6975
R8698 a_n17351_68.n31 a_n17351_68.t24 17.6975
R8699 a_n17351_68.n24 a_n17351_68.t24 17.6975
R8700 a_n17351_68.n32 a_n17351_68.t29 17.6975
R8701 a_n17351_68.n23 a_n17351_68.t29 17.6975
R8702 a_n17351_68.n33 a_n17351_68.t22 17.6975
R8703 a_n17351_68.n22 a_n17351_68.t22 17.6975
R8704 a_n17351_68.n34 a_n17351_68.t26 17.6975
R8705 a_n17351_68.n21 a_n17351_68.t26 17.6975
R8706 a_n17351_68.n35 a_n17351_68.t10 17.6975
R8707 a_n17351_68.n20 a_n17351_68.t10 17.6975
R8708 a_n17351_68.n36 a_n17351_68.t25 17.6975
R8709 a_n17351_68.n19 a_n17351_68.t25 17.6975
R8710 a_n17351_68.t2 a_n17351_68.n1 17.6975
R8711 a_n17351_68.n18 a_n17351_68.t2 17.6975
R8712 a_n17351_68.n2 a_n17351_68.t28 17.6975
R8713 a_n17351_68.n17 a_n17351_68.t28 17.6975
R8714 a_n17351_68.n3 a_n17351_68.t38 17.6975
R8715 a_n17351_68.n16 a_n17351_68.t38 17.6975
R8716 a_n17351_68.n4 a_n17351_68.t20 17.6975
R8717 a_n17351_68.n15 a_n17351_68.t20 17.6975
R8718 a_n17351_68.n5 a_n17351_68.t32 17.6975
R8719 a_n17351_68.n14 a_n17351_68.t32 17.6975
R8720 a_n17351_68.n6 a_n17351_68.t13 17.6975
R8721 a_n17351_68.n13 a_n17351_68.t13 17.6975
R8722 a_n17351_68.n7 a_n17351_68.t30 17.6975
R8723 a_n17351_68.n12 a_n17351_68.t30 17.6975
R8724 a_n17351_68.n8 a_n17351_68.t23 17.6975
R8725 a_n17351_68.n11 a_n17351_68.t23 17.6975
R8726 a_n17351_68.n9 a_n17351_68.t36 17.6975
R8727 a_n17351_68.n10 a_n17351_68.t36 17.6975
R8728 a_n17351_68.n9 a_n17351_68.n8 15.513
R8729 a_n17351_68.n8 a_n17351_68.n7 15.513
R8730 a_n17351_68.n7 a_n17351_68.n6 15.513
R8731 a_n17351_68.n6 a_n17351_68.n5 15.513
R8732 a_n17351_68.n5 a_n17351_68.n4 15.513
R8733 a_n17351_68.n4 a_n17351_68.n3 15.513
R8734 a_n17351_68.n3 a_n17351_68.n2 15.513
R8735 a_n17351_68.n2 a_n17351_68.n1 15.513
R8736 a_n17351_68.n36 a_n17351_68.n35 15.513
R8737 a_n17351_68.n35 a_n17351_68.n34 15.513
R8738 a_n17351_68.n34 a_n17351_68.n33 15.513
R8739 a_n17351_68.n33 a_n17351_68.n32 15.513
R8740 a_n17351_68.n32 a_n17351_68.n31 15.513
R8741 a_n17351_68.n31 a_n17351_68.n30 15.513
R8742 a_n17351_68.n30 a_n17351_68.n29 15.513
R8743 a_n17351_68.n29 a_n17351_68.n28 15.513
R8744 a_n17351_68.n46 a_n17351_68.n45 15.513
R8745 a_n17351_68.n45 a_n17351_68.n44 15.513
R8746 a_n17351_68.n44 a_n17351_68.n43 15.513
R8747 a_n17351_68.n43 a_n17351_68.n42 15.513
R8748 a_n17351_68.n42 a_n17351_68.n41 15.513
R8749 a_n17351_68.n41 a_n17351_68.n40 15.513
R8750 a_n17351_68.n40 a_n17351_68.n39 15.513
R8751 a_n17351_68.n39 a_n17351_68.n38 15.513
R8752 a_n17351_68.n73 a_n17351_68.n72 15.513
R8753 a_n17351_68.n72 a_n17351_68.n71 15.513
R8754 a_n17351_68.n71 a_n17351_68.n70 15.513
R8755 a_n17351_68.n70 a_n17351_68.n69 15.513
R8756 a_n17351_68.n69 a_n17351_68.n68 15.513
R8757 a_n17351_68.n68 a_n17351_68.n67 15.513
R8758 a_n17351_68.n67 a_n17351_68.n66 15.513
R8759 a_n17351_68.n66 a_n17351_68.n65 15.513
R8760 a_n17351_68.n75 a_n17351_68.t0 14.2059
R8761 a_n17351_68.n37 a_n17351_68.n1 7.75675
R8762 a_n17351_68.n37 a_n17351_68.n36 7.75675
R8763 a_n17351_68.n74 a_n17351_68.n38 7.75675
R8764 a_n17351_68.n74 a_n17351_68.n73 7.75675
R8765 a_n17351_68.t1 a_n17351_68.n75 4.23734
R8766 a_n17351_68.n0 a_n17351_68.n37 0.633736
R8767 a_n17351_68.n0 a_n17351_68.n74 0.59343
R8768 a_n17351_68.n0 a_n17351_68.n75 2.39173
R8769 a_22203_n358.n5 a_22203_n358.t15 31.6987
R8770 a_22203_n358.n6 a_22203_n358.t17 18.6885
R8771 a_22203_n358.n7 a_22203_n358.t14 18.6885
R8772 a_22203_n358.n5 a_22203_n358.t18 18.6885
R8773 a_22203_n358.n10 a_22203_n358.t16 13.907
R8774 a_22203_n358.n9 a_22203_n358.t12 13.8462
R8775 a_22203_n358.n11 a_22203_n358.t20 13.8462
R8776 a_22203_n358.n9 a_22203_n358.t9 12.1185
R8777 a_22203_n358.n11 a_22203_n358.t19 12.1185
R8778 a_22203_n358.n10 a_22203_n358.t8 12.0455
R8779 a_22203_n358.n6 a_22203_n358.t10 11.1938
R8780 a_22203_n358.n7 a_22203_n358.t13 11.1938
R8781 a_22203_n358.n5 a_22203_n358.t11 11.1938
R8782 a_22203_n358.n1 a_22203_n358.n9 10.6383
R8783 a_22203_n358.n7 a_22203_n358.n6 10.5449
R8784 a_22203_n358.n1 a_22203_n358.n11 10.2813
R8785 a_22203_n358.n1 a_22203_n358.n10 10.2813
R8786 a_22203_n358.n0 a_22203_n358.n4 7.33746
R8787 a_22203_n358.n8 a_22203_n358.n5 6.48939
R8788 a_22203_n358.n0 a_22203_n358.n3 6.46093
R8789 a_22203_n358.n12 a_22203_n358.n0 6.01368
R8790 a_22203_n358.n0 a_22203_n358.n2 5.4118
R8791 a_22203_n358.n8 a_22203_n358.n7 4.05606
R8792 a_22203_n358.n4 a_22203_n358.t0 3.6005
R8793 a_22203_n358.n4 a_22203_n358.t3 3.6005
R8794 a_22203_n358.n3 a_22203_n358.t1 3.6005
R8795 a_22203_n358.n3 a_22203_n358.t2 3.6005
R8796 a_22203_n358.n0 a_22203_n358.n1 2.59067
R8797 a_22203_n358.n0 a_22203_n358.n8 2.22925
R8798 a_22203_n358.n2 a_22203_n358.t4 2.06607
R8799 a_22203_n358.n12 a_22203_n358.t6 2.06607
R8800 a_22203_n358.n2 a_22203_n358.t5 1.4923
R8801 a_22203_n358.t7 a_22203_n358.n12 1.4923
R8802 a_n4208_n141.n2 a_n4208_n141.t4 26.5147
R8803 a_n4208_n141.n1 a_n4208_n141.t3 25.076
R8804 a_n4208_n141.n1 a_n4208_n141.t6 25.076
R8805 a_n4208_n141.n3 a_n4208_n141.t7 25.076
R8806 a_n4208_n141.n3 a_n4208_n141.t8 25.076
R8807 a_n4208_n141.n2 a_n4208_n141.t5 25.076
R8808 a_n4208_n141.n0 a_n4208_n141.t0 23.009
R8809 a_n4208_n141.n0 a_n4208_n141.t1 12.3005
R8810 a_n4208_n141.t2 a_n4208_n141.n1 11.2556
R8811 a_n4208_n141.n1 a_n4208_n141.n0 3.08843
R8812 a_n4208_n141.n1 a_n4208_n141.n3 2.8778
R8813 a_n4208_n141.n3 a_n4208_n141.n2 2.8778
R8814 a_n8471_219.n1 a_n8471_219.t6 31.1854
R8815 a_n8471_219.n0 a_n8471_219.t8 30.4809
R8816 a_n8471_219.n0 a_n8471_219.t7 29.7468
R8817 a_n8471_219.n0 a_n8471_219.t5 29.7468
R8818 a_n8471_219.n2 a_n8471_219.t10 29.7468
R8819 a_n8471_219.n2 a_n8471_219.t11 29.7468
R8820 a_n8471_219.n1 a_n8471_219.t9 29.7468
R8821 a_n8471_219.n3 a_n8471_219.t3 28.2414
R8822 a_n8471_219.n0 a_n8471_219.t2 11.7439
R8823 a_n8471_219.n3 a_n8471_219.t4 8.52921
R8824 a_n8471_219.t0 a_n8471_219.n4 4.50971
R8825 a_n8471_219.n4 a_n8471_219.t1 4.38259
R8826 a_n8471_219.n4 a_n8471_219.n0 3.32162
R8827 a_n8471_219.n0 a_n8471_219.n2 2.8778
R8828 a_n8471_219.n2 a_n8471_219.n1 2.8778
R8829 a_n8471_219.n0 a_n8471_219.n3 2.4541
R8830 PLL_REF_CLK PLL_REF_CLK.n0 20.7258
R8831 PLL_REF_CLK.n0 PLL_REF_CLK.t1 17.3015
R8832 PLL_REF_CLK.n0 PLL_REF_CLK.t0 10.6463
R8833 a_23620_8319.n0 a_23620_8319.t5 56.5589
R8834 a_23620_8319.n1 a_23620_8319.t4 54.6195
R8835 a_23620_8319.n1 a_23620_8319.t3 54.3444
R8836 a_23620_8319.n0 a_23620_8319.t6 54.3444
R8837 a_23620_8319.n3 a_23620_8319.n2 7.32981
R8838 a_23620_8319.n3 a_23620_8319.n1 3.5139
R8839 a_23620_8319.t1 a_23620_8319.n3 1.76266
R8840 a_23620_8319.n2 a_23620_8319.t0 1.6385
R8841 a_23620_8319.n2 a_23620_8319.t2 1.6385
R8842 a_23620_8319.n1 a_23620_8319.n0 1.3316
R8843 a_n8537_n1530.n2 a_n8537_n1530.t13 48.7058
R8844 a_n8537_n1530.n10 a_n8537_n1530.t14 47.5611
R8845 a_n8537_n1530.t6 a_n8537_n1530.n11 47.5611
R8846 a_n8537_n1530.n7 a_n8537_n1530.t5 46.602
R8847 a_n8537_n1530.n6 a_n8537_n1530.t9 46.602
R8848 a_n8537_n1530.n5 a_n8537_n1530.t7 46.602
R8849 a_n8537_n1530.n4 a_n8537_n1530.t12 46.602
R8850 a_n8537_n1530.n3 a_n8537_n1530.t10 46.602
R8851 a_n8537_n1530.n2 a_n8537_n1530.t15 46.602
R8852 a_n8537_n1530.n0 a_n8537_n1530.n13 37.0921
R8853 a_n8537_n1530.t14 a_n8537_n1530.n9 33.9289
R8854 a_n8537_n1530.n12 a_n8537_n1530.t6 33.9289
R8855 a_n8537_n1530.n12 a_n8537_n1530.t11 28.7581
R8856 a_n8537_n1530.n11 a_n8537_n1530.t11 28.7581
R8857 a_n8537_n1530.t4 a_n8537_n1530.n9 28.7581
R8858 a_n8537_n1530.n10 a_n8537_n1530.t4 28.7581
R8859 a_n8537_n1530.n11 a_n8537_n1530.n10 18.8035
R8860 a_n8537_n1530.n17 a_n8537_n1530.t0 6.3005
R8861 a_n8537_n1530.n17 a_n8537_n1530.n16 4.85375
R8862 a_n8537_n1530.n15 a_n8537_n1530.n14 4.5005
R8863 a_n8537_n1530.n1 a_n8537_n1530.n0 1.83275
R8864 a_n8537_n1530.n13 a_n8537_n1530.n9 2.58592
R8865 a_n8537_n1530.n13 a_n8537_n1530.n12 2.58592
R8866 a_n8537_n1530.t2 a_n8537_n1530.n17 2.56843
R8867 a_n8537_n1530.t0 a_n8537_n1530.t3 1.6385
R8868 a_n8537_n1530.n16 a_n8537_n1530.n8 1.51412
R8869 a_n8537_n1530.n3 a_n8537_n1530.n2 1.00625
R8870 a_n8537_n1530.t1 a_n8537_n1530.t2 0.813
R8871 a_n8537_n1530.n7 a_n8537_n1530.n6 0.62375
R8872 a_n8537_n1530.n4 a_n8537_n1530.n3 0.57425
R8873 a_n8537_n1530.n6 a_n8537_n1530.n5 0.57425
R8874 a_n8537_n1530.n5 a_n8537_n1530.n4 0.25475
R8875 a_n8537_n1530.n14 a_n8537_n1530.n8 0.233801
R8876 a_n8537_n1530.n8 a_n8537_n1530.n7 0.169297
R8877 a_n8537_n1530.n15 a_n8537_n1530.n0 0.15575
R8878 a_n8537_n1530.n14 a_n8537_n1530.n1 0.148629
R8879 a_n8537_n1530.n16 a_n8537_n1530.n15 0.11975
R8880 a_n8537_n1530.n1 a_n8537_n1530.t8 46.6222
R8881 a_22115_253.n2 a_22115_253.t5 121.874
R8882 a_22115_253.t5 a_22115_253.t7 61.5152
R8883 a_22115_253.n0 a_22115_253.t4 52.378
R8884 a_22115_253.n0 a_22115_253.t3 17.7152
R8885 a_22115_253.n1 a_22115_253.t0 11.1158
R8886 a_22115_253.n1 a_22115_253.n2 9.95623
R8887 a_22115_253.n1 a_22115_253.n0 8.37615
R8888 a_22115_253.t1 a_22115_253.n1 8.02846
R8889 a_22115_253.n0 a_22115_253.t6 7.36133
R8890 a_22115_253.n2 a_22115_253.t2 6.7165
R8891 a_n8537_93.t4 a_n8537_93.n4 47.5611
R8892 a_n8537_93.n3 a_n8537_93.t12 47.5611
R8893 a_n8537_93.n0 a_n8537_93.n6 36.4925
R8894 a_n8537_93.n5 a_n8537_93.t4 33.9289
R8895 a_n8537_93.t12 a_n8537_93.n2 33.9289
R8896 a_n8537_93.n1 a_n8537_93.t3 31.0687
R8897 a_n8537_93.n0 a_n8537_93.t1 29.4084
R8898 a_n8537_93.n0 a_n8537_93.t14 29.3475
R8899 a_n8537_93.n0 a_n8537_93.t10 29.3475
R8900 a_n8537_93.n0 a_n8537_93.t5 29.3475
R8901 a_n8537_93.n0 a_n8537_93.t8 29.3475
R8902 a_n8537_93.n1 a_n8537_93.t6 29.3475
R8903 a_n8537_93.n1 a_n8537_93.t9 29.3475
R8904 a_n8537_93.n1 a_n8537_93.t7 29.3475
R8905 a_n8537_93.t11 a_n8537_93.n2 28.7581
R8906 a_n8537_93.n3 a_n8537_93.t11 28.7581
R8907 a_n8537_93.n5 a_n8537_93.t13 28.7581
R8908 a_n8537_93.n4 a_n8537_93.t13 28.7581
R8909 a_n8537_93.n4 a_n8537_93.n3 18.8035
R8910 a_n8537_93.n0 a_n8537_93.t2 10.616
R8911 a_n8537_93.t0 a_n8537_93.n0 4.49193
R8912 a_n8537_93.n0 a_n8537_93.n1 3.41375
R8913 a_n8537_93.n6 a_n8537_93.n2 2.58592
R8914 a_n8537_93.n6 a_n8537_93.n5 2.58592
R8915 a_21394_11355.n6 a_21394_11355.t21 50.888
R8916 a_21394_11355.n7 a_21394_11355.t19 50.888
R8917 a_21394_11355.n8 a_21394_11355.t29 50.888
R8918 a_21394_11355.n9 a_21394_11355.t23 50.888
R8919 a_21394_11355.n10 a_21394_11355.t18 50.888
R8920 a_21394_11355.n11 a_21394_11355.t24 50.888
R8921 a_21394_11355.n12 a_21394_11355.t20 50.888
R8922 a_21394_11355.n13 a_21394_11355.t22 50.888
R8923 a_21394_11355.n6 a_21394_11355.t6 50.888
R8924 a_21394_11355.n7 a_21394_11355.t10 50.888
R8925 a_21394_11355.n8 a_21394_11355.t14 50.888
R8926 a_21394_11355.n9 a_21394_11355.t2 50.888
R8927 a_21394_11355.n10 a_21394_11355.t12 50.888
R8928 a_21394_11355.n11 a_21394_11355.t16 50.888
R8929 a_21394_11355.n12 a_21394_11355.t8 50.888
R8930 a_21394_11355.n13 a_21394_11355.t4 50.888
R8931 a_21394_11355.n16 a_21394_11355.t25 29.0305
R8932 a_21394_11355.n15 a_21394_11355.t27 29.0305
R8933 a_21394_11355.n19 a_21394_11355.t28 28.988
R8934 a_21394_11355.n17 a_21394_11355.t26 28.988
R8935 a_21394_11355.n21 a_21394_11355.n20 2.2505
R8936 a_21394_11355.n18 a_21394_11355.n14 2.2505
R8937 a_21394_11355.n1 a_21394_11355.n13 2.05375
R8938 a_21394_11355.n2 a_21394_11355.n5 1.9899
R8939 a_21394_11355.n0 a_21394_11355.n23 1.54264
R8940 a_21394_11355.n1 a_21394_11355.n24 1.51597
R8941 a_21394_11355.n1 a_21394_11355.n4 1.51597
R8942 a_21394_11355.n25 a_21394_11355.n1 1.51457
R8943 a_21394_11355.n16 a_21394_11355.n14 1.16575
R8944 a_21394_11355.n21 a_21394_11355.n15 1.16575
R8945 a_21394_11355.n3 a_21394_11355.n22 0.770928
R8946 a_21394_11355.n1 a_21394_11355.n2 0.0230833
R8947 a_21394_11355.n23 a_21394_11355.t11 0.3255
R8948 a_21394_11355.n23 a_21394_11355.t7 0.3255
R8949 a_21394_11355.n24 a_21394_11355.t3 0.3255
R8950 a_21394_11355.n24 a_21394_11355.t15 0.3255
R8951 a_21394_11355.n4 a_21394_11355.t5 0.3255
R8952 a_21394_11355.n4 a_21394_11355.t9 0.3255
R8953 a_21394_11355.t17 a_21394_11355.n25 0.3255
R8954 a_21394_11355.n25 a_21394_11355.t13 0.3255
R8955 a_21394_11355.n5 a_21394_11355.t0 0.293
R8956 a_21394_11355.n5 a_21394_11355.t1 0.293
R8957 a_21394_11355.n20 a_21394_11355.n18 0.04025
R8958 a_21394_11355.n17 a_21394_11355.n16 0.039655
R8959 a_21394_11355.n19 a_21394_11355.n15 0.039655
R8960 a_21394_11355.n13 a_21394_11355.n12 0.0352143
R8961 a_21394_11355.n12 a_21394_11355.n11 0.0352143
R8962 a_21394_11355.n11 a_21394_11355.n10 0.0352143
R8963 a_21394_11355.n10 a_21394_11355.n9 0.0352143
R8964 a_21394_11355.n8 a_21394_11355.n7 0.0352143
R8965 a_21394_11355.n7 a_21394_11355.n6 0.0352143
R8966 a_21394_11355.n9 a_21394_11355.n8 0.0352143
R8967 a_21394_11355.n18 a_21394_11355.n17 0.021125
R8968 a_21394_11355.n20 a_21394_11355.n19 0.021125
R8969 a_21394_11355.n22 a_21394_11355.n14 0.020375
R8970 a_21394_11355.n22 a_21394_11355.n21 0.020375
R8971 a_21394_11355.n3 a_21394_11355.n2 0.0692465
R8972 a_21394_11355.n3 a_21394_11355.n0 0.147139
R8973 a_21394_11355.n1 a_21394_11355.n0 0.08297
R8974 a_21506_13215.n2 a_21506_13215.t10 51.0134
R8975 a_21506_13215.n2 a_21506_13215.t11 50.7576
R8976 a_21506_13215.n0 a_21506_13215.n1 1.90384
R8977 a_21506_13215.n7 a_21506_13215.n5 1.55709
R8978 a_21506_13215.n7 a_21506_13215.n6 1.51597
R8979 a_21506_13215.n4 a_21506_13215.n3 1.51597
R8980 a_21506_13215.n9 a_21506_13215.n8 1.51457
R8981 a_21506_13215.n0 a_21506_13215.n2 2.67807
R8982 a_21506_13215.n5 a_21506_13215.t8 0.3255
R8983 a_21506_13215.n5 a_21506_13215.t6 0.3255
R8984 a_21506_13215.n6 a_21506_13215.t4 0.3255
R8985 a_21506_13215.n6 a_21506_13215.t2 0.3255
R8986 a_21506_13215.n3 a_21506_13215.t5 0.3255
R8987 a_21506_13215.n3 a_21506_13215.t7 0.3255
R8988 a_21506_13215.n9 a_21506_13215.t3 0.3255
R8989 a_21506_13215.t9 a_21506_13215.n9 0.3255
R8990 a_21506_13215.n1 a_21506_13215.t1 0.293
R8991 a_21506_13215.n1 a_21506_13215.t0 0.293
R8992 a_21506_13215.n8 a_21506_13215.n4 0.0406869
R8993 a_21506_13215.n8 a_21506_13215.n7 0.0402196
R8994 a_21506_13215.n4 a_21506_13215.n0 0.171403
R8995 a_22941_7733.n0 a_22941_7733.t5 42.2199
R8996 a_22941_7733.n1 a_22941_7733.t0 40.4081
R8997 a_22941_7733.n0 a_22941_7733.t6 40.4081
R8998 a_22941_7733.n0 a_22941_7733.t4 40.4081
R8999 a_22941_7733.n0 a_22941_7733.t3 40.4081
R9000 a_22941_7733.t2 a_22941_7733.n1 7.4853
R9001 a_22941_7733.n1 a_22941_7733.t1 5.40883
R9002 a_22941_7733.n1 a_22941_7733.n0 2.96695
R9003 a_22115_1610.n2 a_22115_1610.t7 121.874
R9004 a_22115_1610.t7 a_22115_1610.t4 61.5152
R9005 a_22115_1610.n0 a_22115_1610.t3 52.378
R9006 a_22115_1610.n0 a_22115_1610.t5 17.7882
R9007 a_22115_1610.n1 a_22115_1610.t0 11.1158
R9008 a_22115_1610.n1 a_22115_1610.n2 9.95623
R9009 a_22115_1610.n1 a_22115_1610.n0 8.37615
R9010 a_22115_1610.t1 a_22115_1610.n1 8.02846
R9011 a_22115_1610.n0 a_22115_1610.t2 7.3005
R9012 a_22115_1610.n2 a_22115_1610.t6 6.7165
R9013 a_22115_n302.n2 a_22115_n302.t7 121.874
R9014 a_22115_n302.t7 a_22115_n302.t4 61.5152
R9015 a_22115_n302.n0 a_22115_n302.t2 52.378
R9016 a_22115_n302.n0 a_22115_n302.t3 17.7882
R9017 a_22115_n302.n1 a_22115_n302.t0 11.1158
R9018 a_22115_n302.n1 a_22115_n302.n2 9.95623
R9019 a_22115_n302.n1 a_22115_n302.n0 8.37615
R9020 a_22115_n302.t1 a_22115_n302.n1 8.02846
R9021 a_22115_n302.n0 a_22115_n302.t6 7.3005
R9022 a_22115_n302.n2 a_22115_n302.t5 6.7165
R9023 a_22388_3950.t0 a_22388_3950.n1 21.2275
R9024 a_22388_3950.n1 a_22388_3950.t5 18.9805
R9025 a_22388_3950.n0 a_22388_3950.t4 17.5205
R9026 a_22388_3950.n0 a_22388_3950.t2 11.5588
R9027 a_22388_3950.n1 a_22388_3950.t3 11.4372
R9028 a_22388_3950.t0 a_22388_3950.t1 8.60523
R9029 a_22388_3950.t0 a_22388_3950.n0 8.27396
C0 a_23347_3522 a_23795_3522 0.012552f
C1 a_22963_1518 a_24090_1243 0.011266f
C2 a_23547_4907 VDD 0.332636f
C3 a_22963_217 a_23455_n345 0.046461f
C4 a_31031_1644 PLL_DISABLE 0.018845f
C5 a_21555_3522 VDD 0.405083f
C6 a_24383_217 VDD 0.520925f
C7 a_21755_4018 a_21855_4398 0.586921f
C8 a_21755_4018 a_27491_1710 0.456773f
C9 a_23455_1567 a_23083_1611 0.107446f
C10 a_22527_1197 a_24090_1243 0.416346f
C11 a_22963_1518 a_24383_1567 0.014406f
C12 a_23099_4907 VDD 0.338717f
C13 a_22963_217 a_22527_n715 0.093423f
C14 a_23883_3430 VDD 0.232629f
C15 a_24090_629 VDD 0.370377f
C16 VDD PLL_CLK_OUT 0.921425f
C17 a_25369_6873 a_23508_2038 0.213175f
C18 a_24891_4907 a_25339_4907 0.013103f
C19 a_23508_2038 a_25334_2082 0.010209f
C20 a_22899_3522 a_23347_3522 0.012552f
C21 a_22527_1197 a_24383_1567 0.023074f
C22 a_22963_1518 a_23083_1611 0.240887f
C23 a_25675_477 a_25587_574 0.285629f
C24 a_22651_4907 VDD 0.337108f
C25 a_23435_3430 VDD 0.205239f
C26 a_31391_1688 PLL_DISABLE 0.019219f
C27 a_23083_261 VDD 0.397896f
C28 a_25369_6873 a_25265_6933 0.136975f
C29 a_22963_1518 a_23455_1567 0.018863f
C30 a_22527_1197 a_23083_1611 0.839895f
C31 a_22203_4907 VDD 0.342721f
C32 a_n2908_8493 a_n2908_7613 0.016713f
C33 a_30943_1688 PLL_DISABLE 0.031524f
C34 a_22987_3430 VDD 0.208767f
C35 a_23455_217 VDD 0.186132f
C36 a_26115_6933 a_26049_6873 0.247434f
C37 a_23691_7733 a_23691_6933 0.022218f
C38 a_24675_7463 a_23508_2038 0.011399f
C39 a_24443_4907 a_24891_4907 0.013103f
C40 a_23883_3430 a_22304_2486 0.026153f
C41 a_22451_3522 a_22899_3522 0.012552f
C42 a_5840_10693 a_5840_9813 0.016713f
C43 a_22527_1197 a_23455_1567 1.16391f
C44 a_21755_4907 VDD 0.396379f
C45 a_27491_1710 PLL_DISABLE 0.106211f
C46 a_22539_3430 VDD 0.212862f
C47 a_22963_217 VDD 0.580508f
C48 a_24675_7463 a_25265_6933 0.090359f
C49 a_24675_7463 a_22864_4398 0.013776f
C50 a_23883_3430 a_23795_3522 0.285629f
C51 a_21755_4018 PLL_DISABLE 0.01221f
C52 a_22527_1197 a_22963_1518 0.280621f
C53 a_5840_8933 a_5840_8053 0.016713f
C54 a_25251_4951 VDD 0.203335f
C55 a_22091_3430 VDD 0.215751f
C56 a_22527_574 VDD 1.1139f
C57 a_24675_7463 a_25095_6933 0.012946f
C58 a_25265_7733 a_26795_7733 0.019086f
C59 a_23995_4907 a_24443_4907 0.013103f
C60 a_22003_3522 a_22451_3522 0.012222f
C61 a_23435_3430 a_23795_3522 0.086905f
C62 a_21667_574 a_21667_n786 0.010569f
C63 a_24803_4951 VDD 0.203482f
C64 a_21643_3430 VDD 0.255373f
C65 a_21667_574 VDD 0.278953f
C66 a_25265_7733 a_26115_6933 1.15373f
C67 a_23508_2038 a_24655_2486 0.057075f
C68 a_23435_3430 a_23347_3522 0.285629f
C69 a_24355_4951 VDD 0.203482f
C70 a_25369_6873 a_26049_6873 1.48855f
C71 a_25369_6873 a_21755_4018 0.19878f
C72 a_23547_4907 a_23995_4907 0.013103f
C73 a_22987_3430 a_23347_3522 0.086905f
C74 a_21555_3522 a_22003_3522 0.012222f
C75 a_n9701_6193 VDD 0.588689f
C76 a_23508_2038 a_24207_2486 0.051499f
C77 a_1220_10693 a_1220_9813 0.016713f
C78 a_21855_1126 a_22963_1518 0.107397f
C79 a_23907_4951 VDD 0.203482f
C80 a_21755_477 VDD 0.377703f
C81 a_25095_7733 a_25265_7733 0.019086f
C82 a_1712_13773 a_1220_13333 0.016789f
C83 a_23508_2038 a_22948_2038 0.542819f
C84 a_22987_3430 a_22899_3522 0.285629f
C85 a_21855_1126 a_22527_1197 0.071077f
C86 a_1220_8933 a_1220_8053 0.016713f
C87 a_23459_4951 VDD 0.203629f
C88 a_24675_7463 a_26049_6873 0.024796f
C89 a_25369_6873 a_26115_6933 0.138982f
C90 a_24675_7463 a_21755_4018 0.08148f
C91 a_25251_4951 a_25339_4907 0.285629f
C92 a_23099_4907 a_23547_4907 0.013103f
C93 a_1220_13773 a_1220_13333 0.016789f
C94 a_22539_3430 a_22899_3522 0.086905f
C95 a_21755_1082 a_25587_1610 0.026006f
C96 a_23011_4951 VDD 0.205777f
C97 a_24090_629 a_24383_217 0.493186f
C98 a_25369_6873 a_25265_7733 0.022799f
C99 a_25251_4951 a_24891_4907 0.087174f
C100 a_18673_2840 a_18489_n1138 0.063905f
C101 a_22539_3430 a_22451_3522 0.285629f
C102 a_22563_4951 VDD 0.208263f
C103 a_n9701_6193 DEBUG 0.073173f
C104 a_24675_7463 a_26115_6933 0.266123f
C105 a_24755_6933 a_25265_7733 0.183758f
C106 a_24803_4951 a_24891_4907 0.285629f
C107 a_22651_4907 a_23099_4907 0.013103f
C108 a_23435_3430 a_23883_3430 0.013276f
C109 a_22091_3430 a_22451_3522 0.086742f
C110 a_23508_2038 a_21755_1082 0.235746f
C111 a_22115_4951 VDD 0.219078f
C112 a_24655_4398 VDD 0.444754f
C113 a_25587_1610 VDD 0.355683f
C114 a_24755_6933 a_25095_7733 0.012025f
C115 a_24675_7463 a_25265_7733 0.180056f
C116 a_24803_4951 a_24443_4907 0.087174f
C117 a_11009_2840 a_14657_n1138 0.058694f
C118 a_22091_3430 a_22003_3522 0.285629f
C119 a_22963_217 a_24383_217 0.015243f
C120 a_23455_217 a_24090_629 0.021118f
C121 a_21667_4951 VDD 0.339057f
C122 a_24207_4398 VDD 0.573638f
C123 a_25675_1518 VDD 0.133852f
C124 a_22203_4907 a_22651_4907 0.013103f
C125 a_24355_4951 a_24443_4907 0.285629f
C126 a_11009_2840 a_10825_n1138 0.046681f
C127 a_5840_14213 a_5840_13333 0.016713f
C128 a_21643_3430 a_22003_3522 0.086742f
C129 a_22987_3430 a_23435_3430 0.013276f
C130 a_1712_11133 a_1712_10253 0.016713f
C131 a_22527_574 a_24383_217 0.023074f
C132 a_23455_217 a_23083_261 0.107446f
C133 a_22963_217 a_24090_629 0.010957f
C134 a_23508_2038 VDD 1.7925f
C135 a_31479_1644 VDD 0.141398f
C136 a_24755_6933 a_25369_6873 0.022154f
C137 a_24355_4951 a_23995_4907 0.087174f
C138 a_7177_2840 a_10825_n1138 0.058694f
C139 a_21643_3430 a_21555_3522 0.285629f
C140 a_24866_11400 a_27414_10401 0.023394f
C141 a_21755_1082 a_24090_1243 0.042898f
C142 a_1712_9373 a_1712_8493 0.016713f
C143 a_22963_217 a_23083_261 0.242122f
C144 a_22527_574 a_24090_629 0.416346f
C145 a_22864_4398 VDD 1.01722f
C146 a_25675_n394 a_25587_n302 0.285629f
C147 a_31031_1644 VDD 0.227358f
C148 a_24675_7463 a_25369_6873 1.05794f
C149 a_21755_4907 a_22203_4907 0.013103f
C150 a_23907_4951 a_23995_4907 0.285629f
C151 a_7177_2840 a_6993_n1138 0.046681f
C152 a_23508_2038 a_22864_2486 0.873597f
C153 a_22539_3430 a_22987_3430 0.013276f
C154 a_21755_1082 a_24383_1567 0.249206f
C155 a_22527_574 a_23083_261 0.839895f
C156 a_22963_217 a_23455_217 0.01975f
C157 a_22948_3950 VDD 0.483198f
C158 a_24675_7463 a_24755_6933 1.50376f
C159 a_23907_4951 a_23547_4907 0.087174f
C160 a_24866_11400 VDD 0.112967f
C161 VDD PLL_FREERUN 9.80733f
C162 a_23508_2038 a_22304_2486 0.132024f
C163 a_22864_4398 a_22864_2486 0.013905f
C164 a_21755_1082 a_23083_1611 0.025834f
C165 a_22527_574 a_23455_217 1.16391f
C166 a_22304_4398 VDD 1.32249f
C167 a_24090_1243 VDD 0.372354f
C168 a_31391_1688 VDD 0.336133f
C169 a_23459_4951 a_23547_4907 0.285629f
C170 a_3345_2840 a_6993_n1138 0.058694f
C171 a_1220_13773 a_1712_13773 0.01254f
C172 a_22091_3430 a_22539_3430 0.013276f
C173 a_n2908_11133 a_n2908_10253 0.016713f
C174 a_21755_1082 a_23455_1567 0.032377f
C175 a_22955_6933 VDD 0.017288f
C176 a_22527_574 a_22963_217 0.307596f
C177 a_24383_1567 VDD 0.523241f
C178 a_30943_1688 VDD 0.365252f
C179 a_23459_4951 a_23099_4907 0.087174f
C180 a_3345_2840 a_3161_n1138 0.046681f
C181 a_22304_4398 a_22864_2486 0.173051f
C182 a_21755_1082 a_22963_1518 0.137044f
C183 a_n2908_9373 a_n2908_8493 0.016713f
C184 a_21855_4398 VDD 0.456781f
C185 a_23083_1611 VDD 0.400846f
C186 a_27491_1710 VDD 0.682158f
C187 a_23011_4951 a_23099_4907 0.285629f
C188 a_24803_4951 a_25251_4951 0.013276f
C189 a_n2908_14213 a_n2908_13333 0.016713f
C190 a_21643_3430 a_22091_3430 0.013276f
C191 a_22304_4398 a_22304_2486 0.01764f
C192 a_5840_11573 a_5840_10693 0.016713f
C193 a_21755_1082 a_22527_1197 0.090966f
C194 a_21855_1126 a_23083_n301 0.227561f
C195 a_26049_6873 VDD 0.526193f
C196 PLL_FREERUN DEBUG 2.62362f
C197 VDD PLL_VCTRL 1.50495f
C198 a_25587_1610 a_25675_477 0.010569f
C199 a_21755_4018 VDD 1.75616f
C200 a_23455_1567 VDD 0.186856f
C201 a_23011_4951 a_22651_4907 0.087174f
C202 a_18477_2840 a_18673_2840 0.106065f
C203 a_n487_2840 a_3161_n1138 0.058694f
C204 a_7177_2840 a_11009_2840 0.971124f
C205 a_26795_7733 VDD 0.02976f
C206 a_18489_n1138 VDD 0.119269f
C207 a_22963_1518 VDD 1.21408f
C208 a_23423_n1258 VDD 1.91928f
C209 a_24355_4951 a_24803_4951 0.013276f
C210 a_22563_4951 a_22651_4907 0.285629f
C211 a_n487_2840 a_n671_n1138 0.046681f
C212 a_21755_4018 a_22864_2486 0.045273f
C213 a_26115_6933 VDD 0.066159f
C214 a_21855_1126 a_22527_n715 0.421686f
C215 a_14657_n1138 VDD 0.119269f
C216 a_22527_1197 VDD 1.11698f
C217 a_21855_n1258 VDD 1.06203f
C218 a_22563_4951 a_22203_4907 0.087174f
C219 a_21755_1082 a_21855_1126 0.77448f
C220 a_25265_7733 VDD 1.11074f
C221 a_21755_477 a_21667_574 0.285629f
C222 a_10825_n1138 VDD 0.119269f
C223 VDD PLL_DISABLE 12.5944f
C224 DEBUG PLL_VCTRL 17.1203f
C225 a_23907_4951 a_24355_4951 0.013276f
C226 a_22115_4951 a_22203_4907 0.285629f
C227 a_3345_2840 a_7177_2840 0.971124f
C228 a_14645_2840 a_11009_2840 0.072091f
C229 a_1220_11573 a_1220_10693 0.016713f
C230 a_22963_1518 a_25587_574 0.023971f
C231 a_25095_7733 VDD 0.02907f
C232 a_31391_1688 PLL_REF_CLK 0.010937f
C233 a_6993_n1138 VDD 0.119269f
C234 a_22115_4951 a_21755_4907 0.087174f
C235 a_25339_4907 a_21755_4018 0.020034f
C236 a_23508_2038 a_23435_3430 0.014853f
C237 a_22304_2486 a_22527_1197 0.010446f
C238 a_24207_2486 a_24655_2486 0.480927f
C239 a_23691_7733 VDD 0.82092f
C240 a_30943_1688 PLL_REF_CLK 0.010937f
C241 a_3161_n1138 VDD 0.119269f
C242 a_24383_n345 a_24090_n669 0.493186f
C243 a_21855_1126 VDD 0.827537f
C244 a_23459_4951 a_23907_4951 0.013276f
C245 a_21667_4951 a_21755_4907 0.285629f
C246 a_10813_2840 a_11009_2840 0.099479f
C247 a_24891_4907 a_21755_4018 0.018929f
C248 a_1712_14653 a_1712_13773 0.016713f
C249 a_25369_6873 VDD 0.86387f
C250 a_27491_1710 PLL_REF_CLK 0.625212f
C251 a_n671_n1138 VDD 0.119269f
C252 a_25587_n302 VDD 0.361795f
C253 a_10813_2840 a_7177_2840 0.072091f
C254 a_24443_4907 a_21755_4018 0.017642f
C255 a_21755_4018 PLL_REF_CLK 0.087887f
C256 a_24755_6933 VDD 1.07973f
C257 a_n8659_n1230 VDD 0.38527f
C258 a_23455_n345 a_24090_n669 0.021118f
C259 a_25675_n394 VDD 0.131378f
C260 a_23011_4951 a_23459_4951 0.013276f
C261 a_23995_4907 a_21755_4018 0.017642f
C262 a_n487_2840 a_3345_2840 0.971124f
C263 a_1220_14653 a_1220_13773 0.016713f
C264 a_22948_3950 a_22987_3430 0.010389f
C265 a_5840_9813 a_5840_8933 0.016713f
C266 a_24675_7463 VDD 1.20178f
C267 a_18673_2840 VDD 0.347176f
C268 a_22527_n715 a_24090_n669 0.416346f
C269 a_23547_4907 a_21755_4018 0.018636f
C270 a_6981_2840 a_7177_2840 0.099479f
C271 a_1220_12453 a_1712_11133 0.016758f
C272 a_22963_1518 a_25675_477 0.010299f
C273 a_11009_2840 VDD 0.629273f
C274 a_22527_n715 a_24383_n345 0.023074f
C275 a_23455_n345 a_23083_n301 0.107446f
C276 a_22563_4951 a_23011_4951 0.013276f
C277 a_23099_4907 a_21755_4018 0.019521f
C278 a_23508_2038 a_25334_3994 0.010314f
C279 PLL_REF_CLK PLL_DISABLE 1.77779f
C280 a_22963_1518 a_24383_217 0.24646f
C281 a_7177_2840 VDD 0.629273f
C282 a_22527_n715 a_23083_n301 0.839895f
C283 a_25587_574 a_25675_n394 0.010569f
C284 a_6981_2840 a_3345_2840 0.072091f
C285 a_22651_4907 a_21755_4018 0.020814f
C286 a_21755_1082 a_22948_2038 0.060492f
C287 a_22963_1518 a_24090_629 0.051285f
C288 a_18477_2840 VDD 0.298308f
C289 a_22527_n715 a_23455_n345 1.16391f
C290 a_24655_2486 VDD 0.443621f
C291 a_24090_n669 VDD 0.371422f
C292 a_22115_4951 a_22563_4951 0.013276f
C293 a_22203_4907 a_21755_4018 0.02231f
C294 a_1220_9813 a_1220_8933 0.016713f
C295 a_22963_1518 a_23083_261 0.045667f
C296 a_3345_2840 VDD 0.629273f
C297 a_24207_2486 VDD 0.57564f
C298 a_24383_n345 VDD 0.524797f
C299 a_24675_7463 a_25339_4907 0.015573f
C300 a_3149_2840 a_3345_2840 0.099479f
C301 a_21755_4907 a_21755_4018 0.010443f
C302 a_n2908_12013 a_n2908_11133 0.016713f
C303 a_22864_2486 a_24655_2486 0.232395f
C304 a_21755_1082 a_21855_2486 0.517726f
C305 a_22963_1518 a_23455_217 0.026991f
C306 a_14645_2840 VDD 0.298285f
C307 PLL_DISABLE PLL_CLK_OUT 2.52613f
C308 a_22948_2038 VDD 0.472672f
C309 a_23083_n301 VDD 0.397859f
C310 a_21667_4951 a_22115_4951 0.013276f
C311 a_25251_4951 a_21755_4018 0.020436f
C312 a_24207_4398 a_24655_4398 0.480927f
C313 a_1220_12453 a_1220_11573 0.024172f
C314 a_22864_2486 a_24207_2486 0.099075f
C315 a_25675_1518 a_25587_1610 0.285629f
C316 a_22963_1518 a_22963_217 0.154909f
C317 a_n487_2840 VDD 0.629273f
C318 a_22963_217 a_23423_n1258 0.016058f
C319 a_23455_n345 VDD 0.186107f
C320 a_3149_2840 a_n487_2840 0.072091f
C321 a_24803_4951 a_21755_4018 0.02016f
C322 a_23508_2038 a_24655_4398 0.05477f
C323 a_22864_2486 a_22948_2038 0.827579f
C324 a_22304_2486 a_24207_2486 0.524f
C325 a_22963_1518 a_22527_574 0.098711f
C326 a_10813_2840 VDD 0.298285f
C327 a_21855_2486 VDD 0.465743f
C328 a_22527_n715 VDD 1.11099f
C329 a_24355_4951 a_21755_4018 0.019809f
C330 a_n683_2840 a_n487_2840 0.099479f
C331 a_1220_14653 a_1712_14653 0.01254f
C332 a_23508_2038 a_24207_4398 0.050704f
C333 a_22864_4398 a_24655_4398 0.224841f
C334 a_22304_2486 a_22948_2038 0.318976f
C335 a_21755_1082 VDD 1.49699f
C336 a_23907_4951 a_21755_4018 0.019809f
C337 a_22864_4398 a_24207_4398 0.097396f
C338 a_27014_14933 a_27814_14933 0.017628f
C339 a_6981_2840 VDD 0.298285f
C340 a_21667_n786 a_21755_n830 0.285629f
C341 a_21755_n830 VDD 0.37735f
C342 a_23459_4951 a_21755_4018 0.020336f
C343 a_22864_4398 a_23508_2038 1.28745f
C344 a_22304_4398 a_24655_4398 0.041108f
C345 a_22304_2486 a_21855_2486 0.051973f
C346 a_1712_10253 a_1712_9373 0.016713f
C347 a_21855_1126 a_22963_217 0.147928f
C348 a_31031_1644 a_31479_1644 0.013276f
C349 a_21667_n786 VDD 0.278953f
C350 a_23011_4951 a_21755_4018 0.020722f
C351 a_22948_3950 a_23508_2038 0.542819f
C352 a_22304_4398 a_24207_4398 0.524441f
C353 a_22304_2486 a_21755_1082 0.029378f
C354 a_21855_1126 a_22527_574 0.075252f
C355 a_3149_2840 VDD 0.298285f
C356 a_22963_217 a_25587_n302 0.024151f
C357 a_22563_4951 a_21755_4018 0.02155f
C358 a_22948_3950 a_22864_4398 0.827579f
C359 a_22304_4398 a_23508_2038 0.290117f
C360 a_n683_2840 VDD 0.298285f
C361 a_22864_2486 VDD 1.0905f
C362 a_31391_1688 a_31479_1644 0.285629f
C363 a_22115_4951 a_21755_4018 0.021129f
C364 a_22304_4398 a_22864_4398 0.79492f
C365 a_24383_217 a_24383_n345 0.01024f
C366 a_31391_1688 a_31031_1644 0.086742f
C367 a_22304_2486 VDD 1.48563f
C368 a_25587_574 VDD 0.222895f
C369 a_24675_7463 a_25251_4951 0.012056f
C370 a_22304_4398 a_22948_3950 0.318865f
C371 a_1220_13333 a_1220_12453 0.041784f
C372 VDD DEBUG 6.47742f
C373 a_n2908_10253 a_n2908_9373 0.016713f
C374 a_23795_3522 VDD 0.340986f
C375 a_30943_1688 a_31031_1644 0.285629f
C376 a_21755_4018 a_23508_2038 0.020593f
C377 a_22304_2486 a_22864_2486 0.77678f
C378 a_25339_4907 VDD 0.337435f
C379 a_23347_3522 VDD 0.332254f
C380 a_26049_6873 a_25265_6933 0.111757f
C381 a_21755_4018 a_22864_4398 0.064811f
C382 a_24383_1567 a_24090_1243 0.493186f
C383 a_24891_4907 VDD 0.333625f
C384 a_22963_217 a_24090_n669 0.05056f
C385 a_22899_3522 VDD 0.336412f
C386 a_30943_1688 a_31391_1688 0.012222f
C387 a_21855_4398 a_22304_4398 0.049604f
C388 a_23795_3522 a_22304_2486 0.019418f
C389 a_22963_217 a_24383_n345 0.266557f
C390 a_24443_4907 VDD 0.331821f
C391 VDD PLL_REF_CLK 1.28796f
C392 a_22451_3522 VDD 0.343186f
C393 PLL_FREERUN PLL_VCTRL 1.34591f
C394 a_26115_6933 a_25265_6933 0.394051f
C395 a_21755_4018 a_22304_4398 0.294635f
C396 a_23347_3522 a_22304_2486 0.011215f
C397 a_23455_1567 a_24090_1243 0.021118f
C398 a_1712_8493 a_1712_7613 0.016713f
C399 a_23995_4907 VDD 0.33177f
C400 a_22963_217 a_23083_n301 0.032472f
C401 a_31479_1644 PLL_DISABLE 0.018672f
C402 a_22003_3522 VDD 0.346078f
C403 a_25675_477 VDD 0.336735f
C404 a_25265_7733 a_25265_6933 0.09437f
C405 PLL_CLK_OUT VSS 3.96787f
C406 PLL_DISABLE VSS 6.736543f
C407 PLL_REF_CLK VSS 1.67389f
C408 PLL_VCTRL VSS 3.841599f
C409 DEBUG VSS 9.152385f
C410 PLL_FREERUN VSS 15.262243f
C411 VDD VSS 0.37829p
C412 a_31479_1644 VSS 0.571591f
C413 a_31031_1644 VSS 0.495269f
C414 a_31391_1688 VSS 0.322948f
C415 a_30943_1688 VSS 0.313069f
C416 a_27491_1710 VSS 0.756683f
C417 a_23423_n1258 VSS 2.97868f
C418 a_21855_n1258 VSS 1.5783f
C419 a_25587_n302 VSS 0.300786f
C420 a_25675_n394 VSS 0.553612f
C421 a_24090_n669 VSS 0.463372f
C422 a_24383_n345 VSS 0.847615f
C423 a_23083_n301 VSS 0.304138f
C424 a_23455_n345 VSS 0.42522f
C425 a_22527_n715 VSS 1.48041f
C426 a_21755_n830 VSS 0.253834f
C427 a_21667_n786 VSS 0.510899f
C428 a_25587_574 VSS 0.503354f
C429 a_25675_477 VSS 0.29293f
C430 a_24383_217 VSS 0.847727f
C431 a_24090_629 VSS 0.46342f
C432 a_23083_261 VSS 0.304138f
C433 a_23455_217 VSS 0.42522f
C434 a_22963_217 VSS 1.30612f
C435 a_22527_574 VSS 1.47988f
C436 a_21667_574 VSS 0.510899f
C437 a_21755_477 VSS 0.255908f
C438 a_25587_1610 VSS 0.301502f
C439 a_25675_1518 VSS 0.561791f
C440 a_24090_1243 VSS 0.468603f
C441 a_24383_1567 VSS 0.851182f
C442 a_23083_1611 VSS 0.30791f
C443 a_23455_1567 VSS 0.425059f
C444 a_22963_1518 VSS 0.66981f
C445 a_22527_1197 VSS 1.48233f
C446 a_21855_1126 VSS 0.731146f
C447 a_24655_2486 VSS 0.49929f
C448 a_24207_2486 VSS 0.52813f
C449 a_22948_2038 VSS 0.653228f
C450 a_21855_2486 VSS 0.487857f
C451 a_21755_1082 VSS 2.34126f
C452 a_22864_2486 VSS 1.26736f
C453 a_22304_2486 VSS 1.62693f
C454 a_23795_3522 VSS 0.291705f
C455 a_23347_3522 VSS 0.285378f
C456 a_22899_3522 VSS 0.286621f
C457 a_22451_3522 VSS 0.288647f
C458 a_22003_3522 VSS 0.288752f
C459 a_21555_3522 VSS 0.292965f
C460 a_23883_3430 VSS 0.496144f
C461 a_23435_3430 VSS 0.476403f
C462 a_22987_3430 VSS 0.478057f
C463 a_22539_3430 VSS 0.482501f
C464 a_22091_3430 VSS 0.482791f
C465 a_21643_3430 VSS 0.49561f
C466 a_24655_4398 VSS 0.501653f
C467 a_24207_4398 VSS 0.525166f
C468 a_23508_2038 VSS 3.2301f
C469 a_22864_4398 VSS 1.30402f
C470 a_22948_3950 VSS 0.663844f
C471 a_22304_4398 VSS 1.59351f
C472 a_21855_4398 VSS 0.486507f
C473 a_21755_4018 VSS 2.81642f
C474 a_18489_n1138 VSS 0.583015f
C475 a_14657_n1138 VSS 0.59026f
C476 a_10825_n1138 VSS 0.59026f
C477 a_6993_n1138 VSS 0.59026f
C478 a_3161_n1138 VSS 0.59026f
C479 a_n671_n1138 VSS 0.59026f
C480 a_n8659_n1230 VSS 2.04194f
C481 a_18673_2840 VSS 1.12107f
C482 a_11009_2840 VSS 3.50221f
C483 a_7177_2840 VSS 3.50221f
C484 a_18477_2840 VSS 0.393424f
C485 a_3345_2840 VSS 3.50221f
C486 a_14645_2840 VSS 0.393424f
C487 a_n487_2840 VSS 3.48363f
C488 a_10813_2840 VSS 0.393424f
C489 a_6981_2840 VSS 0.393424f
C490 a_3149_2840 VSS 0.393424f
C491 a_n683_2840 VSS 0.393424f
C492 a_25339_4907 VSS 0.44212f
C493 a_24891_4907 VSS 0.284703f
C494 a_24443_4907 VSS 0.284815f
C495 a_23995_4907 VSS 0.284088f
C496 a_23547_4907 VSS 0.284758f
C497 a_23099_4907 VSS 0.285892f
C498 a_22651_4907 VSS 0.283647f
C499 a_22203_4907 VSS 0.28405f
C500 a_21755_4907 VSS 0.294904f
C501 a_25251_4951 VSS 0.502807f
C502 a_24803_4951 VSS 0.487275f
C503 a_24355_4951 VSS 0.489361f
C504 a_23907_4951 VSS 0.486164f
C505 a_23459_4951 VSS 0.487236f
C506 a_23011_4951 VSS 0.486282f
C507 a_22563_4951 VSS 0.48952f
C508 a_22115_4951 VSS 0.486149f
C509 a_21667_4951 VSS 0.52688f
C510 a_26795_6933 VSS 0.012152f
C511 a_25265_6933 VSS 0.65977f
C512 a_23691_6933 VSS 0.682074f
C513 a_22955_6933 VSS 0.677414f
C514 a_21891_6933 VSS 0.606695f
C515 a_26049_6873 VSS 1.2196f
C516 a_26115_6933 VSS 0.152057f
C517 a_25265_7733 VSS 0.166494f
C518 a_23691_7733 VSS 0.055944f
C519 a_25369_6873 VSS 4.66053f
C520 a_24755_6933 VSS 0.642077f
C521 a_24675_7463 VSS 2.77221f
C522 a_n9701_6193 VSS 2.79685f
C523 a_16431_6193 VSS 0.790553f
C524 a_1712_7613 VSS 0.768303f
C525 a_n2908_7613 VSS 0.821503f
C526 a_5840_8053 VSS 0.667177f
C527 a_1220_8053 VSS 0.755702f
C528 a_1712_8493 VSS 0.738449f
C529 a_n2908_8493 VSS 0.80006f
C530 a_5840_8933 VSS 0.666596f
C531 a_1220_8933 VSS 0.73827f
C532 a_1712_9373 VSS 0.738245f
C533 a_n2908_9373 VSS 0.798803f
C534 a_27814_14933 VSS 0.674688f
C535 a_27414_10401 VSS 0.658975f
C536 a_27014_14933 VSS 0.669913f
C537 a_5840_9813 VSS 0.666585f
C538 a_1220_9813 VSS 0.738245f
C539 a_1712_10253 VSS 0.738245f
C540 a_n2908_10253 VSS 0.800006f
C541 a_5840_10693 VSS 0.666585f
C542 a_1220_10693 VSS 0.738245f
C543 a_1712_11133 VSS 0.741641f
C544 a_n2908_11133 VSS 0.798351f
C545 a_5840_11573 VSS 0.677754f
C546 a_1220_11573 VSS 0.755665f
C547 a_1220_12453 VSS 0.933081f
C548 a_n2908_12013 VSS 0.809581f
C549 a_24866_11400 VSS 3.02217f
C550 a_1220_13333 VSS 0.921533f
C551 a_5840_13333 VSS 0.677754f
C552 a_n2908_13333 VSS 0.808528f
C553 a_1712_13773 VSS 0.741641f
C554 a_1220_13773 VSS 0.741701f
C555 a_5840_14213 VSS 0.666585f
C556 a_n2908_14213 VSS 0.799661f
C557 a_1712_14653 VSS 0.75376f
C558 a_1220_14653 VSS 0.755212f
C559 a_22388_3950.t0 VSS 1.25053f
C560 a_22388_3950.t1 VSS 0.048467f
C561 a_22388_3950.t4 VSS 0.077986f
C562 a_22388_3950.t2 VSS 0.042413f
C563 a_22388_3950.n0 VSS 0.079885f
C564 a_22388_3950.t5 VSS 0.078379f
C565 a_22388_3950.t3 VSS 0.060967f
C566 a_22388_3950.n1 VSS 0.46137f
C567 a_22115_n302.t6 VSS 0.043151f
C568 a_22115_n302.n0 VSS 0.221428f
C569 a_22115_n302.n1 VSS 0.803219f
C570 a_22115_n302.t2 VSS 0.144509f
C571 a_22115_n302.t3 VSS 0.127487f
C572 a_22115_n302.t0 VSS 0.047684f
C573 a_22115_n302.t5 VSS 0.020325f
C574 a_22115_n302.t4 VSS 0.127787f
C575 a_22115_n302.t7 VSS 0.401653f
C576 a_22115_n302.n2 VSS 0.257957f
C577 a_22115_n302.t1 VSS 0.1048f
C578 a_22115_1610.t2 VSS 0.041275f
C579 a_22115_1610.n0 VSS 0.211801f
C580 a_22115_1610.n1 VSS 0.768297f
C581 a_22115_1610.t3 VSS 0.138226f
C582 a_22115_1610.t5 VSS 0.121944f
C583 a_22115_1610.t0 VSS 0.045611f
C584 a_22115_1610.t6 VSS 0.019441f
C585 a_22115_1610.t4 VSS 0.122231f
C586 a_22115_1610.t7 VSS 0.38419f
C587 a_22115_1610.n2 VSS 0.246741f
C588 a_22115_1610.t1 VSS 0.100244f
C589 a_22941_7733.t2 VSS 0.178922f
C590 a_22941_7733.n0 VSS 1.87028f
C591 a_22941_7733.n1 VSS 0.91684f
C592 a_22941_7733.t5 VSS 0.157433f
C593 a_22941_7733.t3 VSS 0.137792f
C594 a_22941_7733.t4 VSS 0.137792f
C595 a_22941_7733.t6 VSS 0.137792f
C596 a_22941_7733.t0 VSS 0.036593f
C597 a_22941_7733.t1 VSS 0.026552f
C598 a_21506_13215.n0 VSS 1.78222f
C599 a_21506_13215.t3 VSS 0.036394f
C600 a_21506_13215.t1 VSS 0.036394f
C601 a_21506_13215.t0 VSS 0.036394f
C602 a_21506_13215.n1 VSS 0.113776f
C603 a_21506_13215.t10 VSS 0.124218f
C604 a_21506_13215.t11 VSS 0.123932f
C605 a_21506_13215.n2 VSS 0.219528f
C606 a_21506_13215.t5 VSS 0.036394f
C607 a_21506_13215.t7 VSS 0.036394f
C608 a_21506_13215.n3 VSS 0.12902f
C609 a_21506_13215.n4 VSS 1.39739f
C610 a_21506_13215.t8 VSS 0.036394f
C611 a_21506_13215.t6 VSS 0.036394f
C612 a_21506_13215.n5 VSS 0.1382f
C613 a_21506_13215.t4 VSS 0.036394f
C614 a_21506_13215.t2 VSS 0.036394f
C615 a_21506_13215.n6 VSS 0.12902f
C616 a_21506_13215.n7 VSS 0.897035f
C617 a_21506_13215.n8 VSS 0.55272f
C618 a_21506_13215.n9 VSS 0.129001f
C619 a_21506_13215.t9 VSS 0.036394f
C620 a_21394_11355.n0 VSS 0.428547f
C621 a_21394_11355.n1 VSS 2.03599f
C622 a_21394_11355.n2 VSS 3.2778f
C623 a_21394_11355.n3 VSS 2.94941f
C624 a_21394_11355.t13 VSS 0.028706f
C625 a_21394_11355.t5 VSS 0.028706f
C626 a_21394_11355.t9 VSS 0.028706f
C627 a_21394_11355.n4 VSS 0.101765f
C628 a_21394_11355.t0 VSS 0.028706f
C629 a_21394_11355.t1 VSS 0.028706f
C630 a_21394_11355.n5 VSS 0.191784f
C631 a_21394_11355.t4 VSS 0.097898f
C632 a_21394_11355.t8 VSS 0.097898f
C633 a_21394_11355.t16 VSS 0.097898f
C634 a_21394_11355.t12 VSS 0.097898f
C635 a_21394_11355.t14 VSS 0.097898f
C636 a_21394_11355.t10 VSS 0.097898f
C637 a_21394_11355.t6 VSS 0.097898f
C638 a_21394_11355.t21 VSS 0.097898f
C639 a_21394_11355.n6 VSS 0.148897f
C640 a_21394_11355.t19 VSS 0.097898f
C641 a_21394_11355.n7 VSS 0.18754f
C642 a_21394_11355.t29 VSS 0.097898f
C643 a_21394_11355.n8 VSS 0.187569f
C644 a_21394_11355.t2 VSS 0.097898f
C645 a_21394_11355.t23 VSS 0.097898f
C646 a_21394_11355.n9 VSS 0.199892f
C647 a_21394_11355.t18 VSS 0.097898f
C648 a_21394_11355.n10 VSS 0.18754f
C649 a_21394_11355.t24 VSS 0.097898f
C650 a_21394_11355.n11 VSS 0.18754f
C651 a_21394_11355.t20 VSS 0.097898f
C652 a_21394_11355.n12 VSS 0.18754f
C653 a_21394_11355.t22 VSS 0.097898f
C654 a_21394_11355.n13 VSS 0.264491f
C655 a_21394_11355.n14 VSS 0.076714f
C656 a_21394_11355.t27 VSS 0.042007f
C657 a_21394_11355.n15 VSS 0.063068f
C658 a_21394_11355.t25 VSS 0.042007f
C659 a_21394_11355.n16 VSS 0.063068f
C660 a_21394_11355.t26 VSS 0.041946f
C661 a_21394_11355.n17 VSS 0.037947f
C662 a_21394_11355.n18 VSS 0.019045f
C663 a_21394_11355.t28 VSS 0.041946f
C664 a_21394_11355.n19 VSS 0.037947f
C665 a_21394_11355.n20 VSS 0.019045f
C666 a_21394_11355.n21 VSS 0.076714f
C667 a_21394_11355.n22 VSS 0.639124f
C668 a_21394_11355.t11 VSS 0.028706f
C669 a_21394_11355.t7 VSS 0.028706f
C670 a_21394_11355.n23 VSS 0.106165f
C671 a_21394_11355.t3 VSS 0.028706f
C672 a_21394_11355.t15 VSS 0.028706f
C673 a_21394_11355.n24 VSS 0.101765f
C674 a_21394_11355.n25 VSS 0.101751f
C675 a_21394_11355.t17 VSS 0.028706f
C676 a_n8537_93.n0 VSS 6.09595f
C677 a_n8537_93.n1 VSS 1.08916f
C678 a_n8537_93.t0 VSS 0.287725f
C679 a_n8537_93.t3 VSS 0.060225f
C680 a_n8537_93.t7 VSS 0.038171f
C681 a_n8537_93.t9 VSS 0.038171f
C682 a_n8537_93.t6 VSS 0.038171f
C683 a_n8537_93.t8 VSS 0.038171f
C684 a_n8537_93.t5 VSS 0.038171f
C685 a_n8537_93.t10 VSS 0.038171f
C686 a_n8537_93.t14 VSS 0.038171f
C687 a_n8537_93.t1 VSS 0.012232f
C688 a_n8537_93.n2 VSS 0.232035f
C689 a_n8537_93.t13 VSS 0.056513f
C690 a_n8537_93.t11 VSS 0.056513f
C691 a_n8537_93.t12 VSS 0.096345f
C692 a_n8537_93.n3 VSS 0.097801f
C693 a_n8537_93.n4 VSS 0.097801f
C694 a_n8537_93.t4 VSS 0.096345f
C695 a_n8537_93.n5 VSS 0.232035f
C696 a_n8537_93.n6 VSS 9.97896f
C697 a_n8537_93.t2 VSS 0.04316f
C698 a_22115_253.t6 VSS 0.042682f
C699 a_22115_253.n0 VSS 0.221505f
C700 a_22115_253.n1 VSS 0.803219f
C701 a_22115_253.t7 VSS 0.127787f
C702 a_22115_253.t5 VSS 0.401653f
C703 a_22115_253.t2 VSS 0.020325f
C704 a_22115_253.n2 VSS 0.257957f
C705 a_22115_253.t4 VSS 0.144509f
C706 a_22115_253.t3 VSS 0.127878f
C707 a_22115_253.t0 VSS 0.047684f
C708 a_22115_253.t1 VSS 0.1048f
C709 a_n8537_n1530.n0 VSS 4.12067f
C710 a_n8537_n1530.n1 VSS 0.157388f
C711 a_n8537_n1530.t2 VSS 0.165534f
C712 a_n8537_n1530.t13 VSS 0.057058f
C713 a_n8537_n1530.t15 VSS 0.043005f
C714 a_n8537_n1530.n2 VSS 0.627589f
C715 a_n8537_n1530.t10 VSS 0.043005f
C716 a_n8537_n1530.n3 VSS 0.17591f
C717 a_n8537_n1530.t12 VSS 0.043005f
C718 a_n8537_n1530.n4 VSS 0.106964f
C719 a_n8537_n1530.t7 VSS 0.043005f
C720 a_n8537_n1530.n5 VSS 0.106964f
C721 a_n8537_n1530.t9 VSS 0.043005f
C722 a_n8537_n1530.n6 VSS 0.140818f
C723 a_n8537_n1530.t5 VSS 0.043005f
C724 a_n8537_n1530.n7 VSS 0.110239f
C725 a_n8537_n1530.n8 VSS 0.030516f
C726 a_n8537_n1530.n9 VSS 0.1818f
C727 a_n8537_n1530.t11 VSS 0.044278f
C728 a_n8537_n1530.t4 VSS 0.044278f
C729 a_n8537_n1530.t14 VSS 0.075487f
C730 a_n8537_n1530.n10 VSS 0.076628f
C731 a_n8537_n1530.n11 VSS 0.076628f
C732 a_n8537_n1530.t6 VSS 0.075487f
C733 a_n8537_n1530.n12 VSS 0.1818f
C734 a_n8537_n1530.n13 VSS 9.222469f
C735 a_n8537_n1530.t8 VSS 0.043067f
C736 a_n8537_n1530.n14 VSS 0.0391f
C737 a_n8537_n1530.n15 VSS 0.021881f
C738 a_n8537_n1530.n16 VSS 0.150424f
C739 a_n8537_n1530.t0 VSS 0.040253f
C740 a_n8537_n1530.t3 VSS 0.013418f
C741 a_n8537_n1530.n17 VSS 0.225262f
C742 a_n8537_n1530.t1 VSS 0.030056f
C743 a_23620_8319.t1 VSS 0.230327f
C744 a_23620_8319.n0 VSS 1.12967f
C745 a_23620_8319.n1 VSS 0.948259f
C746 a_23620_8319.t0 VSS 0.02864f
C747 a_23620_8319.t2 VSS 0.02864f
C748 a_23620_8319.n2 VSS 0.085133f
C749 a_23620_8319.t5 VSS 0.160449f
C750 a_23620_8319.t6 VSS 0.141303f
C751 a_23620_8319.t3 VSS 0.141303f
C752 a_23620_8319.t4 VSS 0.142193f
C753 a_23620_8319.n3 VSS 0.564088f
C754 a_n8471_219.n0 VSS 4.02225f
C755 a_n8471_219.n1 VSS 1.52386f
C756 a_n8471_219.n2 VSS 1.96436f
C757 a_n8471_219.n3 VSS 0.450257f
C758 a_n8471_219.t1 VSS 0.050494f
C759 a_n8471_219.t0 VSS 0.052129f
C760 a_n8471_219.t4 VSS 0.017122f
C761 a_n8471_219.t3 VSS 0.010371f
C762 a_n8471_219.t8 VSS 0.016824f
C763 a_n8471_219.t6 VSS 0.040735f
C764 a_n8471_219.t9 VSS 0.014537f
C765 a_n8471_219.t11 VSS 0.014537f
C766 a_n8471_219.t10 VSS 0.014537f
C767 a_n8471_219.t5 VSS 0.014537f
C768 a_n8471_219.t7 VSS 0.014537f
C769 a_n8471_219.t2 VSS 0.031516f
C770 a_n8471_219.n4 VSS 0.6474f
C771 a_n4208_n141.n0 VSS 0.168853f
C772 a_n4208_n141.n1 VSS 2.09118f
C773 a_n4208_n141.n2 VSS 0.918953f
C774 a_n4208_n141.n3 VSS 1.17828f
C775 a_n4208_n141.t4 VSS 0.026767f
C776 a_n4208_n141.t2 VSS 0.069682f
C777 a_22203_n358.n0 VSS 0.603745f
C778 a_22203_n358.n1 VSS 1.31566f
C779 a_22203_n358.t6 VSS 0.018938f
C780 a_22203_n358.t4 VSS 0.018938f
C781 a_22203_n358.t5 VSS 0.013677f
C782 a_22203_n358.n2 VSS 0.032956f
C783 a_22203_n358.n3 VSS 0.010391f
C784 a_22203_n358.n4 VSS 0.014693f
C785 a_22203_n358.t15 VSS 0.054532f
C786 a_22203_n358.t18 VSS 0.035955f
C787 a_22203_n358.t11 VSS 0.020179f
C788 a_22203_n358.n5 VSS 0.096198f
C789 a_22203_n358.t17 VSS 0.035955f
C790 a_22203_n358.t10 VSS 0.020179f
C791 a_22203_n358.n6 VSS 0.062148f
C792 a_22203_n358.t14 VSS 0.035955f
C793 a_22203_n358.t13 VSS 0.020179f
C794 a_22203_n358.n7 VSS 0.065252f
C795 a_22203_n358.n8 VSS 0.041506f
C796 a_22203_n358.t12 VSS 0.025088f
C797 a_22203_n358.t9 VSS 0.026733f
C798 a_22203_n358.n9 VSS 0.058633f
C799 a_22203_n358.t8 VSS 0.026841f
C800 a_22203_n358.t16 VSS 0.024974f
C801 a_22203_n358.n10 VSS 0.048595f
C802 a_22203_n358.t20 VSS 0.025088f
C803 a_22203_n358.t19 VSS 0.026733f
C804 a_22203_n358.n11 VSS 0.048589f
C805 a_22203_n358.n12 VSS 0.037604f
C806 a_22203_n358.t7 VSS 0.013677f
C807 a_n17351_68.n0 VSS 9.27113f
C808 a_n17351_68.t0 VSS 0.056057f
C809 a_n17351_68.n1 VSS 0.032323f
C810 a_n17351_68.t25 VSS 0.02205f
C811 a_n17351_68.t10 VSS 0.02205f
C812 a_n17351_68.t26 VSS 0.02205f
C813 a_n17351_68.t22 VSS 0.02205f
C814 a_n17351_68.t29 VSS 0.02205f
C815 a_n17351_68.t24 VSS 0.02205f
C816 a_n17351_68.t31 VSS 0.02205f
C817 a_n17351_68.t18 VSS 0.02205f
C818 a_n17351_68.t33 VSS 0.02205f
C819 a_n17351_68.t2 VSS 0.02205f
C820 a_n17351_68.t28 VSS 0.02205f
C821 a_n17351_68.t38 VSS 0.02205f
C822 a_n17351_68.t20 VSS 0.02205f
C823 a_n17351_68.t32 VSS 0.02205f
C824 a_n17351_68.t13 VSS 0.02205f
C825 a_n17351_68.t30 VSS 0.02205f
C826 a_n17351_68.t23 VSS 0.02205f
C827 a_n17351_68.t36 VSS 0.02205f
C828 a_n17351_68.n2 VSS 0.039423f
C829 a_n17351_68.n3 VSS 0.039423f
C830 a_n17351_68.n4 VSS 0.039423f
C831 a_n17351_68.n5 VSS 0.039423f
C832 a_n17351_68.n6 VSS 0.039423f
C833 a_n17351_68.n7 VSS 0.039423f
C834 a_n17351_68.n8 VSS 0.039423f
C835 a_n17351_68.n9 VSS 0.055801f
C836 a_n17351_68.t35 VSS 0.050464f
C837 a_n17351_68.n10 VSS 0.047683f
C838 a_n17351_68.n11 VSS 0.034453f
C839 a_n17351_68.n12 VSS 0.034453f
C840 a_n17351_68.n13 VSS 0.034453f
C841 a_n17351_68.n14 VSS 0.034453f
C842 a_n17351_68.n15 VSS 0.034453f
C843 a_n17351_68.n16 VSS 0.034453f
C844 a_n17351_68.n17 VSS 0.034453f
C845 a_n17351_68.n18 VSS 0.034453f
C846 a_n17351_68.n19 VSS 0.034453f
C847 a_n17351_68.n20 VSS 0.034453f
C848 a_n17351_68.n21 VSS 0.034453f
C849 a_n17351_68.n22 VSS 0.034453f
C850 a_n17351_68.n23 VSS 0.034453f
C851 a_n17351_68.n24 VSS 0.034453f
C852 a_n17351_68.n25 VSS 0.034453f
C853 a_n17351_68.n26 VSS 0.034453f
C854 a_n17351_68.n27 VSS 0.047683f
C855 a_n17351_68.t27 VSS 0.050464f
C856 a_n17351_68.n28 VSS 0.055801f
C857 a_n17351_68.n29 VSS 0.039423f
C858 a_n17351_68.n30 VSS 0.039423f
C859 a_n17351_68.n31 VSS 0.039423f
C860 a_n17351_68.n32 VSS 0.039423f
C861 a_n17351_68.n33 VSS 0.039423f
C862 a_n17351_68.n34 VSS 0.039423f
C863 a_n17351_68.n35 VSS 0.039423f
C864 a_n17351_68.n36 VSS 0.032323f
C865 a_n17351_68.n37 VSS 0.588605f
C866 a_n17351_68.n38 VSS 0.046104f
C867 a_n17351_68.t5 VSS 0.049612f
C868 a_n17351_68.t4 VSS 0.049612f
C869 a_n17351_68.t41 VSS 0.049612f
C870 a_n17351_68.t19 VSS 0.049612f
C871 a_n17351_68.t17 VSS 0.049612f
C872 a_n17351_68.t16 VSS 0.049612f
C873 a_n17351_68.t11 VSS 0.049612f
C874 a_n17351_68.t7 VSS 0.049612f
C875 a_n17351_68.t6 VSS 0.049612f
C876 a_n17351_68.t9 VSS 0.049612f
C877 a_n17351_68.t14 VSS 0.049612f
C878 a_n17351_68.t15 VSS 0.049612f
C879 a_n17351_68.t37 VSS 0.049612f
C880 a_n17351_68.t39 VSS 0.049612f
C881 a_n17351_68.t40 VSS 0.049612f
C882 a_n17351_68.t3 VSS 0.049612f
C883 a_n17351_68.t8 VSS 0.049612f
C884 a_n17351_68.t12 VSS 0.049612f
C885 a_n17351_68.n39 VSS 0.053204f
C886 a_n17351_68.n40 VSS 0.053204f
C887 a_n17351_68.n41 VSS 0.053204f
C888 a_n17351_68.n42 VSS 0.053204f
C889 a_n17351_68.n43 VSS 0.053204f
C890 a_n17351_68.n44 VSS 0.053204f
C891 a_n17351_68.n45 VSS 0.053204f
C892 a_n17351_68.n46 VSS 0.08524f
C893 a_n17351_68.t34 VSS 0.075266f
C894 a_n17351_68.n47 VSS 0.076129f
C895 a_n17351_68.n48 VSS 0.048234f
C896 a_n17351_68.n49 VSS 0.048234f
C897 a_n17351_68.n50 VSS 0.048234f
C898 a_n17351_68.n51 VSS 0.048234f
C899 a_n17351_68.n52 VSS 0.048234f
C900 a_n17351_68.n53 VSS 0.048234f
C901 a_n17351_68.n54 VSS 0.048234f
C902 a_n17351_68.n55 VSS 0.048234f
C903 a_n17351_68.n56 VSS 0.048234f
C904 a_n17351_68.n57 VSS 0.048234f
C905 a_n17351_68.n58 VSS 0.048234f
C906 a_n17351_68.n59 VSS 0.048234f
C907 a_n17351_68.n60 VSS 0.048234f
C908 a_n17351_68.n61 VSS 0.048234f
C909 a_n17351_68.n62 VSS 0.048234f
C910 a_n17351_68.n63 VSS 0.048234f
C911 a_n17351_68.n64 VSS 0.076129f
C912 a_n17351_68.t21 VSS 0.075266f
C913 a_n17351_68.n65 VSS 0.08524f
C914 a_n17351_68.n66 VSS 0.053204f
C915 a_n17351_68.n67 VSS 0.053204f
C916 a_n17351_68.n68 VSS 0.053204f
C917 a_n17351_68.n69 VSS 0.053204f
C918 a_n17351_68.n70 VSS 0.053204f
C919 a_n17351_68.n71 VSS 0.053204f
C920 a_n17351_68.n72 VSS 0.053204f
C921 a_n17351_68.n73 VSS 0.046104f
C922 a_n17351_68.n74 VSS 0.241226f
C923 a_n17351_68.n75 VSS 0.660994f
C924 a_n17351_68.t1 VSS 0.234287f
C925 a_n558_2704.n0 VSS 0.767275f
C926 a_n558_2704.n1 VSS 0.10249f
C927 a_n558_2704.n2 VSS 1.15531f
C928 a_n558_2704.t1 VSS 0.011378f
C929 a_n558_2704.n3 VSS 1.09908f
C930 a_n558_2704.t0 VSS 0.017613f
C931 a_n15085_2072.n1 VSS 0.043242f
C932 a_n15085_2072.n4 VSS 0.037357f
C933 a_n15085_2072.n6 VSS 10.506599f
C934 a_n15085_2072.n9 VSS 0.015756f
C935 a_n15085_2072.n11 VSS 0.019809f
C936 a_n15085_2072.n12 VSS 3.06204f
C937 a_n15085_2072.n14 VSS 0.010493f
C938 a_n15085_2072.n23 VSS 0.029924f
C939 a_n15085_2072.n26 VSS 0.03094f
C940 a_n15085_2072.n27 VSS 0.03094f
C941 a_n15085_2072.n29 VSS 0.030827f
C942 a_n15085_2072.n30 VSS 0.030789f
C943 a_n15085_2072.n31 VSS 0.030051f
C944 a_n15085_2072.n32 VSS 0.030051f
C945 a_n15085_2072.n34 VSS 0.029924f
C946 a_n15085_2072.t20 VSS 0.012567f
C947 a_n15085_2072.t48 VSS 0.262536f
C948 a_n15085_2072.t49 VSS 0.262536f
C949 a_n15085_2072.t47 VSS 0.262536f
C950 a_n15085_2072.t41 VSS 0.262536f
C951 a_n15085_2072.t42 VSS 0.262536f
C952 a_n15085_2072.t43 VSS 0.262536f
C953 a_n15085_2072.t44 VSS 0.262536f
C954 a_n15085_2072.t50 VSS 0.262536f
C955 a_n15085_2072.t45 VSS 0.262536f
C956 a_n15085_2072.t46 VSS 0.262536f
C957 PLL_DISABLE.n0 VSS 0.104716f
C958 PLL_DISABLE.t21 VSS 0.112683f
C959 PLL_DISABLE.t2 VSS 0.112683f
C960 PLL_DISABLE.t15 VSS 0.112683f
C961 PLL_DISABLE.t14 VSS 0.112683f
C962 PLL_DISABLE.t34 VSS 0.112683f
C963 PLL_DISABLE.t11 VSS 0.112683f
C964 PLL_DISABLE.t4 VSS 0.112683f
C965 PLL_DISABLE.t17 VSS 0.112683f
C966 PLL_DISABLE.t1 VSS 0.112683f
C967 PLL_DISABLE.t30 VSS 0.112683f
C968 PLL_DISABLE.t12 VSS 0.112683f
C969 PLL_DISABLE.t36 VSS 0.112683f
C970 PLL_DISABLE.t26 VSS 0.112683f
C971 PLL_DISABLE.t0 VSS 0.112683f
C972 PLL_DISABLE.t16 VSS 0.112683f
C973 PLL_DISABLE.t3 VSS 0.112683f
C974 PLL_DISABLE.t9 VSS 0.112683f
C975 PLL_DISABLE.t31 VSS 0.112683f
C976 PLL_DISABLE.n1 VSS 0.12084f
C977 PLL_DISABLE.n2 VSS 0.12084f
C978 PLL_DISABLE.n3 VSS 0.12084f
C979 PLL_DISABLE.n4 VSS 0.12084f
C980 PLL_DISABLE.n5 VSS 0.12084f
C981 PLL_DISABLE.n6 VSS 0.12084f
C982 PLL_DISABLE.n7 VSS 0.12084f
C983 PLL_DISABLE.n8 VSS 0.193604f
C984 PLL_DISABLE.t7 VSS 0.17095f
C985 PLL_DISABLE.n9 VSS 0.172911f
C986 PLL_DISABLE.n10 VSS 0.109553f
C987 PLL_DISABLE.n11 VSS 0.109553f
C988 PLL_DISABLE.n12 VSS 0.109553f
C989 PLL_DISABLE.n13 VSS 0.109553f
C990 PLL_DISABLE.n14 VSS 0.109553f
C991 PLL_DISABLE.n15 VSS 0.109553f
C992 PLL_DISABLE.n16 VSS 0.109553f
C993 PLL_DISABLE.n17 VSS 0.109553f
C994 PLL_DISABLE.n18 VSS 0.109553f
C995 PLL_DISABLE.n19 VSS 0.109553f
C996 PLL_DISABLE.n20 VSS 0.109553f
C997 PLL_DISABLE.n21 VSS 0.109553f
C998 PLL_DISABLE.n22 VSS 0.109553f
C999 PLL_DISABLE.n23 VSS 0.109553f
C1000 PLL_DISABLE.n24 VSS 0.109553f
C1001 PLL_DISABLE.n25 VSS 0.109553f
C1002 PLL_DISABLE.n26 VSS 0.172911f
C1003 PLL_DISABLE.t19 VSS 0.17095f
C1004 PLL_DISABLE.n27 VSS 0.193604f
C1005 PLL_DISABLE.n28 VSS 0.12084f
C1006 PLL_DISABLE.n29 VSS 0.12084f
C1007 PLL_DISABLE.n30 VSS 0.12084f
C1008 PLL_DISABLE.n31 VSS 0.12084f
C1009 PLL_DISABLE.n32 VSS 0.12084f
C1010 PLL_DISABLE.n33 VSS 0.12084f
C1011 PLL_DISABLE.n34 VSS 0.12084f
C1012 PLL_DISABLE.n35 VSS 0.104716f
C1013 PLL_DISABLE.n36 VSS 4.20208f
C1014 PLL_DISABLE.t5 VSS 0.039814f
C1015 PLL_DISABLE.t37 VSS 0.040419f
C1016 PLL_DISABLE.n37 VSS 0.138474f
C1017 PLL_DISABLE.n38 VSS 1.6969f
C1018 PLL_DISABLE.n39 VSS 0.518544f
C1019 PLL_DISABLE.t20 VSS 0.087706f
C1020 PLL_DISABLE.t23 VSS 0.085935f
C1021 PLL_DISABLE.n40 VSS 0.138154f
C1022 PLL_DISABLE.t10 VSS 0.087706f
C1023 PLL_DISABLE.t29 VSS 0.085935f
C1024 PLL_DISABLE.n41 VSS 0.145154f
C1025 PLL_DISABLE.t13 VSS 0.087706f
C1026 PLL_DISABLE.t33 VSS 0.085935f
C1027 PLL_DISABLE.n42 VSS 0.138154f
C1028 PLL_DISABLE.t25 VSS 0.087706f
C1029 PLL_DISABLE.t32 VSS 0.085935f
C1030 PLL_DISABLE.n43 VSS 0.141739f
C1031 PLL_DISABLE.n44 VSS 0.296935f
C1032 PLL_DISABLE.t6 VSS 0.087706f
C1033 PLL_DISABLE.t24 VSS 0.085935f
C1034 PLL_DISABLE.n45 VSS 0.152324f
C1035 PLL_DISABLE.t28 VSS 0.087706f
C1036 PLL_DISABLE.t35 VSS 0.085935f
C1037 PLL_DISABLE.n46 VSS 0.15591f
C1038 PLL_DISABLE.t8 VSS 0.087706f
C1039 PLL_DISABLE.t27 VSS 0.085935f
C1040 PLL_DISABLE.n47 VSS 0.15591f
C1041 PLL_DISABLE.t18 VSS 0.087706f
C1042 PLL_DISABLE.t22 VSS 0.085935f
C1043 PLL_DISABLE.n48 VSS 0.14891f
C1044 PLL_DISABLE.n49 VSS 0.301872f
C1045 PLL_DISABLE.n50 VSS 1.29015f
C1046 DEBUG.t80 VSS 0.218204f
C1047 DEBUG.t45 VSS 0.458682f
C1048 DEBUG.t14 VSS 0.121237f
C1049 DEBUG.t78 VSS 0.071456f
C1050 DEBUG.t68 VSS 0.071456f
C1051 DEBUG.n0 VSS 0.348853f
C1052 DEBUG.t13 VSS 0.023819f
C1053 DEBUG.t23 VSS 0.023819f
C1054 DEBUG.n1 VSS 0.068817f
C1055 DEBUG.t63 VSS 0.071456f
C1056 DEBUG.t48 VSS 0.071456f
C1057 DEBUG.n2 VSS 0.348853f
C1058 DEBUG.t10 VSS 0.023819f
C1059 DEBUG.t20 VSS 0.023819f
C1060 DEBUG.n3 VSS 0.068817f
C1061 DEBUG.t47 VSS 0.071456f
C1062 DEBUG.t42 VSS 0.071456f
C1063 DEBUG.n4 VSS 0.348853f
C1064 DEBUG.t17 VSS 0.023819f
C1065 DEBUG.t24 VSS 0.023819f
C1066 DEBUG.n5 VSS 0.068817f
C1067 DEBUG.t75 VSS 0.071456f
C1068 DEBUG.t74 VSS 0.071456f
C1069 DEBUG.n6 VSS 0.348853f
C1070 DEBUG.t18 VSS 0.023819f
C1071 DEBUG.t12 VSS 0.023819f
C1072 DEBUG.n7 VSS 0.068817f
C1073 DEBUG.t69 VSS 0.071456f
C1074 DEBUG.t52 VSS 0.071456f
C1075 DEBUG.n8 VSS 0.348853f
C1076 DEBUG.t22 VSS 0.023819f
C1077 DEBUG.t9 VSS 0.023819f
C1078 DEBUG.n9 VSS 0.068817f
C1079 DEBUG.t64 VSS 0.071456f
C1080 DEBUG.t61 VSS 0.071456f
C1081 DEBUG.n10 VSS 0.348853f
C1082 DEBUG.t6 VSS 0.023819f
C1083 DEBUG.t15 VSS 0.023819f
C1084 DEBUG.n11 VSS 0.068817f
C1085 DEBUG.t57 VSS 0.071456f
C1086 DEBUG.t55 VSS 0.071456f
C1087 DEBUG.n12 VSS 0.348853f
C1088 DEBUG.t7 VSS 0.023819f
C1089 DEBUG.t16 VSS 0.023819f
C1090 DEBUG.n13 VSS 0.068817f
C1091 DEBUG.t76 VSS 0.071456f
C1092 DEBUG.t77 VSS 0.071456f
C1093 DEBUG.n14 VSS 0.348853f
C1094 DEBUG.t11 VSS 0.023819f
C1095 DEBUG.t21 VSS 0.023819f
C1096 DEBUG.n15 VSS 0.068817f
C1097 DEBUG.t54 VSS 0.071456f
C1098 DEBUG.t53 VSS 0.071456f
C1099 DEBUG.n16 VSS 0.348853f
C1100 DEBUG.t8 VSS 0.023819f
C1101 DEBUG.t25 VSS 0.023819f
C1102 DEBUG.n17 VSS 0.068817f
C1103 DEBUG.t59 VSS 0.458682f
C1104 DEBUG.t19 VSS 0.121237f
C1105 DEBUG.n18 VSS 0.996133f
C1106 DEBUG.n19 VSS 0.991652f
C1107 DEBUG.n20 VSS 0.976995f
C1108 DEBUG.n21 VSS 0.976995f
C1109 DEBUG.n22 VSS 0.976995f
C1110 DEBUG.n23 VSS 0.976995f
C1111 DEBUG.n24 VSS 0.976995f
C1112 DEBUG.n25 VSS 0.976995f
C1113 DEBUG.n26 VSS 0.976995f
C1114 DEBUG.n27 VSS 0.991652f
C1115 DEBUG.n28 VSS 2.81029f
C1116 DEBUG.t5 VSS 0.458682f
C1117 DEBUG.t40 VSS 0.121237f
C1118 DEBUG.t4 VSS 0.071456f
C1119 DEBUG.t33 VSS 0.071456f
C1120 DEBUG.n29 VSS 0.348853f
C1121 DEBUG.t41 VSS 0.023819f
C1122 DEBUG.t49 VSS 0.023819f
C1123 DEBUG.n30 VSS 0.068817f
C1124 DEBUG.t26 VSS 0.071456f
C1125 DEBUG.t0 VSS 0.071456f
C1126 DEBUG.n31 VSS 0.348853f
C1127 DEBUG.t72 VSS 0.023819f
C1128 DEBUG.t79 VSS 0.023819f
C1129 DEBUG.n32 VSS 0.068817f
C1130 DEBUG.t38 VSS 0.071456f
C1131 DEBUG.t35 VSS 0.071456f
C1132 DEBUG.n33 VSS 0.348853f
C1133 DEBUG.t43 VSS 0.023819f
C1134 DEBUG.t58 VSS 0.023819f
C1135 DEBUG.n34 VSS 0.068817f
C1136 DEBUG.t3 VSS 0.071456f
C1137 DEBUG.t28 VSS 0.071456f
C1138 DEBUG.n35 VSS 0.348853f
C1139 DEBUG.t46 VSS 0.023819f
C1140 DEBUG.t67 VSS 0.023819f
C1141 DEBUG.n36 VSS 0.068817f
C1142 DEBUG.t2 VSS 0.071456f
C1143 DEBUG.t31 VSS 0.071456f
C1144 DEBUG.n37 VSS 0.348853f
C1145 DEBUG.t62 VSS 0.023819f
C1146 DEBUG.t51 VSS 0.023819f
C1147 DEBUG.n38 VSS 0.068817f
C1148 DEBUG.t1 VSS 0.071456f
C1149 DEBUG.t30 VSS 0.071456f
C1150 DEBUG.n39 VSS 0.348853f
C1151 DEBUG.t70 VSS 0.023819f
C1152 DEBUG.t65 VSS 0.023819f
C1153 DEBUG.n40 VSS 0.068817f
C1154 DEBUG.t34 VSS 0.071456f
C1155 DEBUG.t27 VSS 0.071456f
C1156 DEBUG.n41 VSS 0.348853f
C1157 DEBUG.t60 VSS 0.023819f
C1158 DEBUG.t71 VSS 0.023819f
C1159 DEBUG.n42 VSS 0.068817f
C1160 DEBUG.t32 VSS 0.071456f
C1161 DEBUG.t39 VSS 0.071456f
C1162 DEBUG.n43 VSS 0.348853f
C1163 DEBUG.t50 VSS 0.023819f
C1164 DEBUG.t73 VSS 0.023819f
C1165 DEBUG.n44 VSS 0.068817f
C1166 DEBUG.t36 VSS 0.071456f
C1167 DEBUG.t37 VSS 0.071456f
C1168 DEBUG.n45 VSS 0.348853f
C1169 DEBUG.t56 VSS 0.023819f
C1170 DEBUG.t44 VSS 0.023819f
C1171 DEBUG.n46 VSS 0.068817f
C1172 DEBUG.t29 VSS 0.458682f
C1173 DEBUG.t66 VSS 0.121237f
C1174 DEBUG.n47 VSS 0.996133f
C1175 DEBUG.n48 VSS 0.991652f
C1176 DEBUG.n49 VSS 0.976995f
C1177 DEBUG.n50 VSS 0.976995f
C1178 DEBUG.n51 VSS 0.976995f
C1179 DEBUG.n52 VSS 0.976995f
C1180 DEBUG.n53 VSS 0.976995f
C1181 DEBUG.n54 VSS 0.976995f
C1182 DEBUG.n55 VSS 0.976995f
C1183 DEBUG.n56 VSS 0.991652f
C1184 DEBUG.n57 VSS 1.17523f
C1185 DEBUG.n58 VSS 6.32273f
C1186 PLL_VCTRL.t21 VSS 0.033703f
C1187 PLL_VCTRL.t39 VSS 0.033703f
C1188 PLL_VCTRL.n0 VSS 0.153157f
C1189 PLL_VCTRL.t2 VSS 0.011234f
C1190 PLL_VCTRL.t19 VSS 0.011234f
C1191 PLL_VCTRL.n1 VSS 0.034669f
C1192 PLL_VCTRL.n2 VSS 1.03707f
C1193 PLL_VCTRL.t33 VSS 0.033703f
C1194 PLL_VCTRL.t31 VSS 0.033703f
C1195 PLL_VCTRL.n3 VSS 0.153157f
C1196 PLL_VCTRL.t7 VSS 0.011234f
C1197 PLL_VCTRL.t10 VSS 0.011234f
C1198 PLL_VCTRL.n4 VSS 0.034669f
C1199 PLL_VCTRL.n5 VSS 1.61901f
C1200 PLL_VCTRL.t23 VSS 0.033703f
C1201 PLL_VCTRL.t22 VSS 0.033703f
C1202 PLL_VCTRL.n6 VSS 0.153157f
C1203 PLL_VCTRL.t16 VSS 0.011234f
C1204 PLL_VCTRL.t13 VSS 0.011234f
C1205 PLL_VCTRL.n7 VSS 0.034669f
C1206 PLL_VCTRL.n8 VSS 1.61901f
C1207 PLL_VCTRL.t20 VSS 0.033703f
C1208 PLL_VCTRL.t36 VSS 0.033703f
C1209 PLL_VCTRL.n9 VSS 0.153157f
C1210 PLL_VCTRL.t14 VSS 0.011234f
C1211 PLL_VCTRL.t0 VSS 0.011234f
C1212 PLL_VCTRL.n10 VSS 0.034669f
C1213 PLL_VCTRL.n11 VSS 1.61901f
C1214 PLL_VCTRL.t35 VSS 0.033703f
C1215 PLL_VCTRL.t34 VSS 0.033703f
C1216 PLL_VCTRL.n12 VSS 0.153157f
C1217 PLL_VCTRL.t18 VSS 0.011234f
C1218 PLL_VCTRL.t6 VSS 0.011234f
C1219 PLL_VCTRL.n13 VSS 0.034669f
C1220 PLL_VCTRL.n14 VSS 1.61901f
C1221 PLL_VCTRL.t24 VSS 0.033703f
C1222 PLL_VCTRL.t32 VSS 0.033703f
C1223 PLL_VCTRL.n15 VSS 0.153157f
C1224 PLL_VCTRL.t5 VSS 0.011234f
C1225 PLL_VCTRL.t8 VSS 0.011234f
C1226 PLL_VCTRL.n16 VSS 0.034669f
C1227 PLL_VCTRL.n17 VSS 1.61901f
C1228 PLL_VCTRL.t30 VSS 0.033703f
C1229 PLL_VCTRL.t28 VSS 0.033703f
C1230 PLL_VCTRL.n18 VSS 0.153157f
C1231 PLL_VCTRL.t3 VSS 0.011234f
C1232 PLL_VCTRL.t9 VSS 0.011234f
C1233 PLL_VCTRL.n19 VSS 0.034669f
C1234 PLL_VCTRL.n20 VSS 1.61901f
C1235 PLL_VCTRL.t27 VSS 0.033703f
C1236 PLL_VCTRL.t37 VSS 0.033703f
C1237 PLL_VCTRL.n21 VSS 0.153157f
C1238 PLL_VCTRL.t12 VSS 0.011234f
C1239 PLL_VCTRL.t11 VSS 0.011234f
C1240 PLL_VCTRL.n22 VSS 0.034669f
C1241 PLL_VCTRL.n23 VSS 1.61901f
C1242 PLL_VCTRL.t38 VSS 0.033703f
C1243 PLL_VCTRL.t26 VSS 0.033703f
C1244 PLL_VCTRL.n24 VSS 0.153157f
C1245 PLL_VCTRL.t17 VSS 0.011234f
C1246 PLL_VCTRL.t4 VSS 0.011234f
C1247 PLL_VCTRL.n25 VSS 0.034669f
C1248 PLL_VCTRL.n26 VSS 1.61901f
C1249 PLL_VCTRL.t25 VSS 0.033703f
C1250 PLL_VCTRL.t29 VSS 0.033703f
C1251 PLL_VCTRL.n27 VSS 0.153157f
C1252 PLL_VCTRL.t15 VSS 0.011234f
C1253 PLL_VCTRL.t1 VSS 0.011234f
C1254 PLL_VCTRL.n28 VSS 0.034669f
C1255 PLL_VCTRL.n29 VSS 1.88002f
C1256 PLL_FREERUN.n0 VSS 0.07358f
C1257 PLL_FREERUN.t37 VSS 0.079178f
C1258 PLL_FREERUN.t23 VSS 0.079178f
C1259 PLL_FREERUN.t40 VSS 0.079178f
C1260 PLL_FREERUN.t30 VSS 0.079178f
C1261 PLL_FREERUN.t4 VSS 0.079178f
C1262 PLL_FREERUN.t34 VSS 0.079178f
C1263 PLL_FREERUN.t7 VSS 0.079178f
C1264 PLL_FREERUN.t25 VSS 0.079178f
C1265 PLL_FREERUN.t11 VSS 0.079178f
C1266 PLL_FREERUN.t18 VSS 0.079178f
C1267 PLL_FREERUN.t3 VSS 0.079178f
C1268 PLL_FREERUN.t15 VSS 0.079178f
C1269 PLL_FREERUN.t27 VSS 0.079178f
C1270 PLL_FREERUN.t9 VSS 0.079178f
C1271 PLL_FREERUN.t24 VSS 0.079178f
C1272 PLL_FREERUN.t5 VSS 0.079178f
C1273 PLL_FREERUN.t32 VSS 0.079178f
C1274 PLL_FREERUN.t14 VSS 0.079178f
C1275 PLL_FREERUN.n1 VSS 0.08491f
C1276 PLL_FREERUN.n2 VSS 0.08491f
C1277 PLL_FREERUN.n3 VSS 0.08491f
C1278 PLL_FREERUN.n4 VSS 0.08491f
C1279 PLL_FREERUN.n5 VSS 0.08491f
C1280 PLL_FREERUN.n6 VSS 0.08491f
C1281 PLL_FREERUN.n7 VSS 0.08491f
C1282 PLL_FREERUN.n8 VSS 0.136038f
C1283 PLL_FREERUN.t13 VSS 0.12012f
C1284 PLL_FREERUN.n9 VSS 0.121498f
C1285 PLL_FREERUN.n10 VSS 0.076979f
C1286 PLL_FREERUN.n11 VSS 0.076979f
C1287 PLL_FREERUN.n12 VSS 0.076979f
C1288 PLL_FREERUN.n13 VSS 0.076979f
C1289 PLL_FREERUN.n14 VSS 0.076979f
C1290 PLL_FREERUN.n15 VSS 0.076979f
C1291 PLL_FREERUN.n16 VSS 0.076979f
C1292 PLL_FREERUN.n17 VSS 0.076979f
C1293 PLL_FREERUN.n18 VSS 0.076979f
C1294 PLL_FREERUN.n19 VSS 0.076979f
C1295 PLL_FREERUN.n20 VSS 0.076979f
C1296 PLL_FREERUN.n21 VSS 0.076979f
C1297 PLL_FREERUN.n22 VSS 0.076979f
C1298 PLL_FREERUN.n23 VSS 0.076979f
C1299 PLL_FREERUN.n24 VSS 0.076979f
C1300 PLL_FREERUN.n25 VSS 0.076979f
C1301 PLL_FREERUN.n26 VSS 0.121498f
C1302 PLL_FREERUN.t1 VSS 0.12012f
C1303 PLL_FREERUN.n27 VSS 0.136038f
C1304 PLL_FREERUN.n28 VSS 0.08491f
C1305 PLL_FREERUN.n29 VSS 0.08491f
C1306 PLL_FREERUN.n30 VSS 0.08491f
C1307 PLL_FREERUN.n31 VSS 0.08491f
C1308 PLL_FREERUN.n32 VSS 0.08491f
C1309 PLL_FREERUN.n33 VSS 0.08491f
C1310 PLL_FREERUN.n34 VSS 0.08491f
C1311 PLL_FREERUN.n35 VSS 0.07358f
C1312 PLL_FREERUN.n36 VSS 2.10553f
C1313 PLL_FREERUN.t38 VSS 0.041918f
C1314 PLL_FREERUN.n37 VSS 1.04593f
C1315 PLL_FREERUN.n38 VSS 0.051586f
C1316 PLL_FREERUN.t33 VSS 0.03519f
C1317 PLL_FREERUN.t41 VSS 0.03519f
C1318 PLL_FREERUN.t21 VSS 0.03519f
C1319 PLL_FREERUN.t39 VSS 0.03519f
C1320 PLL_FREERUN.t20 VSS 0.03519f
C1321 PLL_FREERUN.t29 VSS 0.03519f
C1322 PLL_FREERUN.t10 VSS 0.03519f
C1323 PLL_FREERUN.t36 VSS 0.03519f
C1324 PLL_FREERUN.t0 VSS 0.03519f
C1325 PLL_FREERUN.t8 VSS 0.03519f
C1326 PLL_FREERUN.t28 VSS 0.03519f
C1327 PLL_FREERUN.t17 VSS 0.03519f
C1328 PLL_FREERUN.t2 VSS 0.03519f
C1329 PLL_FREERUN.t19 VSS 0.03519f
C1330 PLL_FREERUN.t12 VSS 0.03519f
C1331 PLL_FREERUN.t31 VSS 0.03519f
C1332 PLL_FREERUN.t6 VSS 0.03519f
C1333 PLL_FREERUN.t26 VSS 0.03519f
C1334 PLL_FREERUN.n39 VSS 0.062916f
C1335 PLL_FREERUN.n40 VSS 0.062916f
C1336 PLL_FREERUN.n41 VSS 0.062916f
C1337 PLL_FREERUN.n42 VSS 0.062916f
C1338 PLL_FREERUN.n43 VSS 0.062916f
C1339 PLL_FREERUN.n44 VSS 0.062916f
C1340 PLL_FREERUN.n45 VSS 0.062916f
C1341 PLL_FREERUN.n46 VSS 0.089056f
C1342 PLL_FREERUN.t22 VSS 0.080537f
C1343 PLL_FREERUN.n47 VSS 0.076099f
C1344 PLL_FREERUN.n48 VSS 0.054985f
C1345 PLL_FREERUN.n49 VSS 0.054985f
C1346 PLL_FREERUN.n50 VSS 0.054985f
C1347 PLL_FREERUN.n51 VSS 0.054985f
C1348 PLL_FREERUN.n52 VSS 0.054985f
C1349 PLL_FREERUN.n53 VSS 0.054985f
C1350 PLL_FREERUN.n54 VSS 0.054985f
C1351 PLL_FREERUN.n55 VSS 0.054985f
C1352 PLL_FREERUN.n56 VSS 0.054985f
C1353 PLL_FREERUN.n57 VSS 0.054985f
C1354 PLL_FREERUN.n58 VSS 0.054985f
C1355 PLL_FREERUN.n59 VSS 0.054985f
C1356 PLL_FREERUN.n60 VSS 0.054985f
C1357 PLL_FREERUN.n61 VSS 0.054985f
C1358 PLL_FREERUN.n62 VSS 0.054985f
C1359 PLL_FREERUN.n63 VSS 0.054985f
C1360 PLL_FREERUN.n64 VSS 0.076099f
C1361 PLL_FREERUN.t16 VSS 0.080537f
C1362 PLL_FREERUN.n65 VSS 0.089056f
C1363 PLL_FREERUN.n66 VSS 0.062916f
C1364 PLL_FREERUN.n67 VSS 0.062916f
C1365 PLL_FREERUN.n68 VSS 0.062916f
C1366 PLL_FREERUN.n69 VSS 0.062916f
C1367 PLL_FREERUN.n70 VSS 0.062916f
C1368 PLL_FREERUN.n71 VSS 0.062916f
C1369 PLL_FREERUN.n72 VSS 0.062916f
C1370 PLL_FREERUN.n73 VSS 0.051586f
C1371 PLL_FREERUN.n74 VSS 2.10446f
C1372 PLL_FREERUN.t35 VSS 0.094642f
C1373 PLL_FREERUN.n75 VSS 1.10052f
C1374 PLL_FREERUN.n76 VSS 0.364432f
C1375 a_22388_2038.t1 VSS 1.25053f
C1376 a_22388_2038.t0 VSS 0.048467f
C1377 a_22388_2038.t5 VSS 0.077986f
C1378 a_22388_2038.t3 VSS 0.042413f
C1379 a_22388_2038.n0 VSS 0.079885f
C1380 a_22388_2038.t2 VSS 0.078379f
C1381 a_22388_2038.t4 VSS 0.060967f
C1382 a_22388_2038.n1 VSS 0.46137f
C1383 a_5840_7613.t0 VSS 26.4671f
C1384 a_5840_7613.t1 VSS 0.032928f
C1385 a_5840_15093.n0 VSS 0.273858f
C1386 a_5840_15093.t9 VSS 29.919199f
C1387 a_5840_15093.n1 VSS 0.158576f
C1388 a_5840_15093.n2 VSS 0.094913f
C1389 a_5840_15093.n3 VSS 0.046236f
C1390 a_5840_15093.n32 VSS 0.021497f
C1391 a_5840_15093.n34 VSS 0.027471f
C1392 a_5840_15093.n35 VSS 0.032271f
C1393 a_5840_15093.n36 VSS 0.012073f
C1394 a_5840_15093.n38 VSS 0.01083f
C1395 a_5840_15093.n52 VSS 0.077048f
C1396 a_5840_15093.n110 VSS 0.013273f
C1397 PLL_CLK_OUT.t31 VSS 0.05541f
C1398 PLL_CLK_OUT.t6 VSS 0.05541f
C1399 PLL_CLK_OUT.n0 VSS 0.404595f
C1400 PLL_CLK_OUT.t32 VSS 0.05541f
C1401 PLL_CLK_OUT.t5 VSS 0.05541f
C1402 PLL_CLK_OUT.n1 VSS 0.404595f
C1403 PLL_CLK_OUT.t29 VSS 0.05541f
C1404 PLL_CLK_OUT.t34 VSS 0.05541f
C1405 PLL_CLK_OUT.n2 VSS 0.404595f
C1406 PLL_CLK_OUT.t2 VSS 0.05541f
C1407 PLL_CLK_OUT.t1 VSS 0.05541f
C1408 PLL_CLK_OUT.n3 VSS 0.404595f
C1409 PLL_CLK_OUT.t39 VSS 0.05541f
C1410 PLL_CLK_OUT.t35 VSS 0.05541f
C1411 PLL_CLK_OUT.n4 VSS 0.404595f
C1412 PLL_CLK_OUT.t8 VSS 0.05541f
C1413 PLL_CLK_OUT.t4 VSS 0.05541f
C1414 PLL_CLK_OUT.n5 VSS 0.404595f
C1415 PLL_CLK_OUT.t37 VSS 0.05541f
C1416 PLL_CLK_OUT.t36 VSS 0.05541f
C1417 PLL_CLK_OUT.n6 VSS 0.404595f
C1418 PLL_CLK_OUT.t0 VSS 0.05541f
C1419 PLL_CLK_OUT.t38 VSS 0.05541f
C1420 PLL_CLK_OUT.n7 VSS 0.404595f
C1421 PLL_CLK_OUT.t33 VSS 0.05541f
C1422 PLL_CLK_OUT.t30 VSS 0.05541f
C1423 PLL_CLK_OUT.n8 VSS 0.404595f
C1424 PLL_CLK_OUT.t3 VSS 0.05541f
C1425 PLL_CLK_OUT.t7 VSS 0.05541f
C1426 PLL_CLK_OUT.n9 VSS 0.404595f
C1427 PLL_CLK_OUT.t13 VSS 0.01847f
C1428 PLL_CLK_OUT.t12 VSS 0.01847f
C1429 PLL_CLK_OUT.n10 VSS 0.056998f
C1430 PLL_CLK_OUT.n11 VSS 0.687802f
C1431 PLL_CLK_OUT.t23 VSS 0.01847f
C1432 PLL_CLK_OUT.t9 VSS 0.01847f
C1433 PLL_CLK_OUT.n12 VSS 0.056998f
C1434 PLL_CLK_OUT.n13 VSS 0.780152f
C1435 PLL_CLK_OUT.t21 VSS 0.01847f
C1436 PLL_CLK_OUT.t26 VSS 0.01847f
C1437 PLL_CLK_OUT.n14 VSS 0.056998f
C1438 PLL_CLK_OUT.n15 VSS 0.780152f
C1439 PLL_CLK_OUT.t28 VSS 0.01847f
C1440 PLL_CLK_OUT.t17 VSS 0.01847f
C1441 PLL_CLK_OUT.n16 VSS 0.056998f
C1442 PLL_CLK_OUT.n17 VSS 0.780152f
C1443 PLL_CLK_OUT.t18 VSS 0.01847f
C1444 PLL_CLK_OUT.t22 VSS 0.01847f
C1445 PLL_CLK_OUT.n18 VSS 0.056998f
C1446 PLL_CLK_OUT.n19 VSS 0.780152f
C1447 PLL_CLK_OUT.t16 VSS 0.01847f
C1448 PLL_CLK_OUT.t19 VSS 0.01847f
C1449 PLL_CLK_OUT.n20 VSS 0.056998f
C1450 PLL_CLK_OUT.n21 VSS 0.780152f
C1451 PLL_CLK_OUT.t11 VSS 0.01847f
C1452 PLL_CLK_OUT.t15 VSS 0.01847f
C1453 PLL_CLK_OUT.n22 VSS 0.056998f
C1454 PLL_CLK_OUT.n23 VSS 0.780152f
C1455 PLL_CLK_OUT.t10 VSS 0.01847f
C1456 PLL_CLK_OUT.t14 VSS 0.01847f
C1457 PLL_CLK_OUT.n24 VSS 0.056998f
C1458 PLL_CLK_OUT.n25 VSS 0.780152f
C1459 PLL_CLK_OUT.t27 VSS 0.01847f
C1460 PLL_CLK_OUT.t24 VSS 0.01847f
C1461 PLL_CLK_OUT.n26 VSS 0.056998f
C1462 PLL_CLK_OUT.n27 VSS 0.780152f
C1463 PLL_CLK_OUT.t25 VSS 0.01847f
C1464 PLL_CLK_OUT.t20 VSS 0.01847f
C1465 PLL_CLK_OUT.n28 VSS 0.056998f
C1466 PLL_CLK_OUT.n29 VSS 2.01444f
C1467 a_27899_438.n0 VSS 2.05379f
C1468 a_27899_438.t3 VSS 0.024107f
C1469 a_27899_438.t9 VSS 0.033969f
C1470 a_27899_438.t10 VSS 0.033979f
C1471 a_27899_438.t12 VSS 0.012498f
C1472 a_27899_438.t5 VSS 0.039632f
C1473 a_27899_438.t6 VSS 0.018274f
C1474 a_27899_438.t0 VSS 0.018274f
C1475 a_27899_438.n1 VSS 0.022026f
C1476 a_27899_438.t23 VSS 0.015026f
C1477 a_27899_438.t19 VSS 0.015026f
C1478 a_27899_438.t13 VSS 0.015026f
C1479 a_27899_438.t24 VSS 0.015026f
C1480 a_27899_438.t20 VSS 0.015026f
C1481 a_27899_438.t15 VSS 0.015026f
C1482 a_27899_438.t18 VSS 0.015026f
C1483 a_27899_438.t32 VSS 0.015026f
C1484 a_27899_438.t28 VSS 0.015026f
C1485 a_27899_438.t22 VSS 0.015026f
C1486 a_27899_438.t25 VSS 0.015026f
C1487 a_27899_438.t26 VSS 0.015026f
C1488 a_27899_438.t30 VSS 0.015026f
C1489 a_27899_438.t27 VSS 0.015026f
C1490 a_27899_438.t31 VSS 0.015026f
C1491 a_27899_438.t17 VSS 0.015026f
C1492 a_27899_438.t14 VSS 0.015026f
C1493 a_27899_438.t21 VSS 0.015026f
C1494 a_27899_438.n2 VSS 0.026864f
C1495 a_27899_438.n3 VSS 0.026864f
C1496 a_27899_438.n4 VSS 0.026864f
C1497 a_27899_438.n5 VSS 0.026864f
C1498 a_27899_438.n6 VSS 0.026864f
C1499 a_27899_438.n7 VSS 0.026864f
C1500 a_27899_438.n8 VSS 0.026864f
C1501 a_27899_438.n9 VSS 0.038025f
C1502 a_27899_438.t16 VSS 0.034388f
C1503 a_27899_438.n10 VSS 0.032493f
C1504 a_27899_438.n11 VSS 0.023477f
C1505 a_27899_438.n12 VSS 0.023477f
C1506 a_27899_438.n13 VSS 0.023477f
C1507 a_27899_438.n14 VSS 0.023477f
C1508 a_27899_438.n15 VSS 0.023477f
C1509 a_27899_438.n16 VSS 0.023477f
C1510 a_27899_438.n17 VSS 0.023477f
C1511 a_27899_438.n18 VSS 0.023477f
C1512 a_27899_438.n19 VSS 0.023477f
C1513 a_27899_438.n20 VSS 0.023477f
C1514 a_27899_438.n21 VSS 0.023477f
C1515 a_27899_438.n22 VSS 0.023477f
C1516 a_27899_438.n23 VSS 0.023477f
C1517 a_27899_438.n24 VSS 0.023477f
C1518 a_27899_438.n25 VSS 0.023477f
C1519 a_27899_438.n26 VSS 0.023477f
C1520 a_27899_438.n27 VSS 0.032493f
C1521 a_27899_438.t29 VSS 0.034388f
C1522 a_27899_438.n28 VSS 0.038025f
C1523 a_27899_438.n29 VSS 0.026864f
C1524 a_27899_438.n30 VSS 0.026864f
C1525 a_27899_438.n31 VSS 0.026864f
C1526 a_27899_438.n32 VSS 0.026864f
C1527 a_27899_438.n33 VSS 0.026864f
C1528 a_27899_438.n34 VSS 0.026864f
C1529 a_27899_438.n35 VSS 0.026864f
C1530 a_27899_438.n36 VSS 0.022026f
C1531 a_27899_438.t7 VSS 0.021399f
C1532 a_27899_438.n37 VSS 0.031259f
C1533 a_27899_438.t1 VSS 0.012498f
C1534 a_24355_n1338.n0 VSS 4.51104f
C1535 a_24355_n1338.n1 VSS 5.21285f
C1536 a_24355_n1338.n2 VSS 0.158565f
C1537 a_24355_n1338.n3 VSS 2.46908f
C1538 a_24355_n1338.t30 VSS 0.02997f
C1539 a_24355_n1338.n4 VSS 0.015495f
C1540 a_24355_n1338.t34 VSS 0.02997f
C1541 a_24355_n1338.t32 VSS 0.02997f
C1542 a_24355_n1338.n5 VSS 0.06069f
C1543 a_24355_n1338.n6 VSS 0.015495f
C1544 a_24355_n1338.t50 VSS 0.094661f
C1545 a_24355_n1338.t15 VSS 0.317616f
C1546 a_24355_n1338.t7 VSS 0.017742f
C1547 a_24355_n1338.t49 VSS 0.017742f
C1548 a_24355_n1338.n7 VSS 0.056271f
C1549 a_24355_n1338.t40 VSS 0.053225f
C1550 a_24355_n1338.t8 VSS 0.053225f
C1551 a_24355_n1338.n8 VSS 0.234884f
C1552 a_24355_n1338.t38 VSS 0.017742f
C1553 a_24355_n1338.t43 VSS 0.017742f
C1554 a_24355_n1338.n9 VSS 0.056271f
C1555 a_24355_n1338.t54 VSS 0.053225f
C1556 a_24355_n1338.t46 VSS 0.053225f
C1557 a_24355_n1338.n10 VSS 0.234884f
C1558 a_24355_n1338.t5 VSS 0.017742f
C1559 a_24355_n1338.t12 VSS 0.017742f
C1560 a_24355_n1338.n11 VSS 0.056271f
C1561 a_24355_n1338.t52 VSS 0.053225f
C1562 a_24355_n1338.t0 VSS 0.053225f
C1563 a_24355_n1338.n12 VSS 0.234884f
C1564 a_24355_n1338.t11 VSS 0.017742f
C1565 a_24355_n1338.t36 VSS 0.017742f
C1566 a_24355_n1338.n13 VSS 0.056271f
C1567 a_24355_n1338.t9 VSS 0.053225f
C1568 a_24355_n1338.t53 VSS 0.053225f
C1569 a_24355_n1338.n14 VSS 0.234884f
C1570 a_24355_n1338.t3 VSS 0.017742f
C1571 a_24355_n1338.t4 VSS 0.017742f
C1572 a_24355_n1338.n15 VSS 0.056271f
C1573 a_24355_n1338.t48 VSS 0.053225f
C1574 a_24355_n1338.t16 VSS 0.053225f
C1575 a_24355_n1338.n16 VSS 0.234884f
C1576 a_24355_n1338.t18 VSS 0.017742f
C1577 a_24355_n1338.t17 VSS 0.017742f
C1578 a_24355_n1338.n17 VSS 0.056271f
C1579 a_24355_n1338.t1 VSS 0.053225f
C1580 a_24355_n1338.t55 VSS 0.053225f
C1581 a_24355_n1338.n18 VSS 0.234884f
C1582 a_24355_n1338.t19 VSS 0.017742f
C1583 a_24355_n1338.t51 VSS 0.017742f
C1584 a_24355_n1338.n19 VSS 0.056271f
C1585 a_24355_n1338.t47 VSS 0.053225f
C1586 a_24355_n1338.t2 VSS 0.053225f
C1587 a_24355_n1338.n20 VSS 0.234884f
C1588 a_24355_n1338.t42 VSS 0.017742f
C1589 a_24355_n1338.t6 VSS 0.017742f
C1590 a_24355_n1338.n21 VSS 0.056271f
C1591 a_24355_n1338.t10 VSS 0.053225f
C1592 a_24355_n1338.t39 VSS 0.053225f
C1593 a_24355_n1338.n22 VSS 0.234884f
C1594 a_24355_n1338.t13 VSS 0.017742f
C1595 a_24355_n1338.t37 VSS 0.017742f
C1596 a_24355_n1338.n23 VSS 0.056271f
C1597 a_24355_n1338.t14 VSS 0.053225f
C1598 a_24355_n1338.t45 VSS 0.053225f
C1599 a_24355_n1338.n24 VSS 0.234884f
C1600 a_24355_n1338.t41 VSS 0.094661f
C1601 a_24355_n1338.t44 VSS 0.317616f
C1602 a_24355_n1338.n25 VSS 0.015495f
C1603 a_24355_n1338.n26 VSS 0.021858f
C1604 a_24355_n1338.t28 VSS 0.02997f
C1605 a_24355_n1338.t33 VSS 0.02997f
C1606 a_24355_n1338.n27 VSS 0.06069f
C1607 a_24355_n1338.t31 VSS 0.02997f
C1608 a_24355_n1338.t29 VSS 0.02997f
C1609 a_24355_n1338.n28 VSS 0.074903f
C1610 a_24355_n1338.n29 VSS 0.06069f
C1611 a_24355_n1338.t35 VSS 0.02997f
C1612 VDD.n0 VSS 0.067687f
C1613 VDD.n1 VSS 0.016922f
C1614 VDD.n2 VSS 0.016922f
C1615 VDD.n3 VSS 0.067687f
C1616 VDD.n4 VSS 0.016922f
C1617 VDD.n5 VSS 0.067687f
C1618 VDD.n6 VSS 0.09287f
C1619 VDD.n7 VSS 0.093133f
C1620 VDD.n8 VSS 0.093133f
C1621 VDD.n9 VSS 0.016922f
C1622 VDD.n10 VSS 0.050826f
C1623 VDD.n11 VSS 0.012852f
C1624 VDD.n12 VSS 0.012852f
C1625 VDD.n13 VSS 0.012852f
C1626 VDD.t38 VSS 0.13974f
C1627 VDD.t262 VSS 0.102581f
C1628 VDD.n14 VSS 0.099117f
C1629 VDD.n15 VSS 0.012852f
C1630 VDD.n16 VSS 0.012852f
C1631 VDD.n17 VSS 0.012852f
C1632 VDD.n18 VSS 0.012852f
C1633 VDD.n20 VSS 0.012852f
C1634 VDD.n21 VSS 0.012852f
C1635 VDD.n23 VSS 0.012852f
C1636 VDD.n24 VSS 0.012852f
C1637 VDD.n26 VSS 0.012852f
C1638 VDD.n27 VSS 0.012852f
C1639 VDD.n29 VSS 0.012852f
C1640 VDD.t142 VSS 0.079814f
C1641 VDD.t363 VSS 0.058618f
C1642 VDD.t270 VSS 0.058618f
C1643 VDD.t280 VSS 0.058618f
C1644 VDD.t336 VSS 0.058618f
C1645 VDD.t285 VSS 0.058618f
C1646 VDD.t87 VSS 0.058618f
C1647 VDD.t359 VSS 0.069347f
C1648 VDD.t19 VSS 0.114095f
C1649 VDD.t21 VSS 0.063328f
C1650 VDD.t145 VSS 0.076674f
C1651 VDD.t284 VSS 0.06673f
C1652 VDD.n30 VSS 0.068762f
C1653 VDD.n31 VSS 0.024027f
C1654 VDD.n32 VSS 0.012852f
C1655 VDD.n33 VSS 0.06796f
C1656 VDD.n34 VSS 0.010415f
C1657 VDD.n35 VSS 0.065158f
C1658 VDD.n36 VSS 0.025429f
C1659 VDD.n38 VSS 0.012852f
C1660 VDD.n39 VSS 0.012852f
C1661 VDD.n40 VSS 0.012852f
C1662 VDD.n41 VSS 0.012852f
C1663 VDD.n42 VSS 0.012852f
C1664 VDD.n43 VSS 0.012852f
C1665 VDD.n44 VSS 0.012791f
C1666 VDD.n45 VSS 0.012852f
C1667 VDD.n46 VSS 0.012852f
C1668 VDD.n47 VSS 0.012852f
C1669 VDD.n48 VSS 0.011094f
C1670 VDD.n49 VSS 0.013394f
C1671 VDD.n51 VSS 0.012852f
C1672 VDD.n52 VSS 0.012852f
C1673 VDD.n53 VSS 0.012852f
C1674 VDD.n54 VSS 0.012852f
C1675 VDD.n55 VSS 0.012549f
C1676 VDD.n58 VSS 0.012852f
C1677 VDD.n59 VSS 0.012852f
C1678 VDD.n60 VSS 0.012852f
C1679 VDD.n61 VSS 0.012852f
C1680 VDD.n62 VSS 0.012852f
C1681 VDD.n65 VSS 0.0117f
C1682 VDD.n66 VSS 0.012852f
C1683 VDD.n67 VSS 0.012852f
C1684 VDD.n68 VSS 0.012852f
C1685 VDD.n69 VSS 0.012852f
C1686 VDD.n72 VSS 0.010245f
C1687 VDD.n73 VSS 0.012852f
C1688 VDD.n74 VSS 0.012852f
C1689 VDD.n75 VSS 0.012852f
C1690 VDD.n76 VSS 0.012852f
C1691 VDD.n77 VSS 0.010488f
C1692 VDD.n78 VSS 0.013416f
C1693 VDD.n80 VSS 0.012852f
C1694 VDD.n81 VSS 0.012852f
C1695 VDD.n82 VSS 0.012852f
C1696 VDD.n84 VSS 0.024028f
C1697 VDD.n85 VSS 0.011154f
C1698 VDD.n86 VSS 0.014068f
C1699 VDD.n88 VSS 0.012852f
C1700 VDD.n89 VSS 0.012852f
C1701 VDD.n90 VSS 0.012852f
C1702 VDD.n91 VSS 0.012852f
C1703 VDD.n92 VSS 0.012852f
C1704 VDD.n94 VSS 0.021372f
C1705 VDD.n95 VSS 0.302029f
C1706 VDD.n96 VSS 0.067687f
C1707 VDD.n97 VSS 0.016922f
C1708 VDD.n98 VSS 0.067687f
C1709 VDD.n99 VSS 0.016922f
C1710 VDD.n100 VSS 0.067687f
C1711 VDD.n101 VSS 0.016922f
C1712 VDD.n102 VSS 0.067687f
C1713 VDD.n103 VSS 0.012851f
C1714 VDD.n104 VSS 0.067687f
C1715 VDD.n106 VSS 0.016922f
C1716 VDD.n107 VSS 0.067687f
C1717 VDD.n108 VSS 0.016922f
C1718 VDD.n109 VSS 0.016922f
C1719 VDD.n110 VSS 0.067687f
C1720 VDD.n111 VSS 0.067687f
C1721 VDD.n112 VSS 0.067687f
C1722 VDD.n113 VSS 0.016922f
C1723 VDD.n114 VSS 0.016922f
C1724 VDD.n115 VSS 0.012532f
C1725 VDD.n116 VSS 0.067687f
C1726 VDD.n117 VSS 0.067687f
C1727 VDD.n118 VSS 0.067687f
C1728 VDD.n119 VSS 0.016922f
C1729 VDD.n120 VSS 0.016922f
C1730 VDD.n121 VSS 0.016922f
C1731 VDD.n122 VSS 0.067687f
C1732 VDD.n123 VSS 0.067687f
C1733 VDD.n124 VSS 0.067687f
C1734 VDD.n125 VSS 0.016922f
C1735 VDD.n126 VSS 0.016922f
C1736 VDD.n127 VSS 0.016922f
C1737 VDD.n128 VSS 0.067687f
C1738 VDD.n129 VSS 0.067687f
C1739 VDD.n130 VSS 0.067687f
C1740 VDD.n131 VSS 0.016922f
C1741 VDD.n132 VSS 0.016922f
C1742 VDD.n133 VSS 0.016922f
C1743 VDD.n134 VSS 0.067687f
C1744 VDD.n135 VSS 0.067687f
C1745 VDD.n136 VSS 0.067687f
C1746 VDD.n137 VSS 0.016922f
C1747 VDD.n138 VSS 0.016922f
C1748 VDD.n139 VSS 0.016922f
C1749 VDD.n140 VSS 0.067687f
C1750 VDD.n141 VSS 0.067687f
C1751 VDD.n142 VSS 0.992578f
C1752 VDD.n143 VSS 0.033418f
C1753 VDD.n144 VSS 0.059499f
C1754 VDD.n145 VSS 0.419585f
C1755 VDD.t279 VSS 0.188689f
C1756 VDD.t122 VSS 0.13638f
C1757 VDD.t282 VSS 0.13638f
C1758 VDD.t114 VSS 0.13638f
C1759 VDD.t268 VSS 0.13638f
C1760 VDD.t327 VSS 0.13638f
C1761 VDD.t89 VSS 0.13638f
C1762 VDD.t63 VSS 0.13638f
C1763 VDD.t366 VSS 0.13638f
C1764 VDD.t338 VSS 0.102285f
C1765 VDD.n146 VSS 0.06819f
C1766 VDD.t144 VSS 0.102285f
C1767 VDD.t113 VSS 0.13638f
C1768 VDD.t362 VSS 0.13638f
C1769 VDD.t361 VSS 0.13638f
C1770 VDD.t62 VSS 0.13638f
C1771 VDD.t365 VSS 0.13638f
C1772 VDD.t283 VSS 0.13638f
C1773 VDD.t269 VSS 0.13638f
C1774 VDD.t112 VSS 0.13638f
C1775 VDD.t141 VSS 0.188689f
C1776 VDD.n147 VSS 0.419585f
C1777 VDD.n148 VSS 0.057546f
C1778 VDD.n149 VSS 0.032942f
C1779 VDD.n150 VSS 7.23992f
C1780 VDD.n151 VSS 0.068627f
C1781 VDD.n152 VSS 1.68476f
C1782 VDD.n153 VSS 0.204207f
C1783 VDD.t255 VSS 0.077475f
C1784 VDD.t254 VSS 0.072269f
C1785 VDD.n159 VSS 0.048695f
C1786 VDD.t157 VSS 0.014711f
C1787 VDD.t212 VSS 0.014711f
C1788 VDD.n161 VSS 0.05179f
C1789 VDD.n162 VSS 0.028927f
C1790 VDD.n167 VSS 0.048695f
C1791 VDD.t214 VSS 0.014711f
C1792 VDD.t245 VSS 0.014711f
C1793 VDD.n169 VSS 0.05179f
C1794 VDD.n170 VSS 0.028927f
C1795 VDD.n175 VSS 0.048695f
C1796 VDD.t174 VSS 0.014711f
C1797 VDD.t257 VSS 0.014711f
C1798 VDD.n177 VSS 0.05179f
C1799 VDD.n178 VSS 0.028927f
C1800 VDD.t253 VSS 0.077984f
C1801 VDD.n184 VSS 0.012099f
C1802 VDD.n186 VSS 0.050672f
C1803 VDD.n187 VSS 0.172582f
C1804 VDD.t252 VSS 0.061763f
C1805 VDD.n188 VSS 0.048695f
C1806 VDD.t173 VSS 0.044194f
C1807 VDD.n189 VSS 0.083886f
C1808 VDD.n201 VSS 0.083886f
C1809 VDD.t256 VSS 0.044194f
C1810 VDD.n202 VSS 0.048695f
C1811 VDD.t213 VSS 0.044194f
C1812 VDD.n203 VSS 0.083886f
C1813 VDD.n215 VSS 0.083886f
C1814 VDD.t244 VSS 0.044194f
C1815 VDD.n216 VSS 0.048695f
C1816 VDD.t156 VSS 0.044194f
C1817 VDD.n217 VSS 0.083886f
C1818 VDD.n230 VSS 0.083886f
C1819 VDD.t211 VSS 0.044194f
C1820 VDD.n231 VSS 0.048695f
C1821 VDD.n232 VSS 0.083886f
C1822 VDD.n235 VSS 0.124948f
C1823 VDD.n236 VSS 0.124605f
C1824 VDD.n238 VSS 0.020742f
C1825 VDD.n239 VSS 0.020464f
C1826 VDD.t275 VSS 0.018109f
C1827 VDD.n240 VSS 0.025135f
C1828 VDD.t82 VSS 0.070455f
C1829 VDD.n241 VSS 0.028468f
C1830 VDD.n242 VSS 0.254273f
C1831 VDD.n243 VSS 0.028468f
C1832 VDD.n244 VSS 0.186579f
C1833 VDD.t353 VSS 0.038983f
C1834 VDD.n245 VSS 0.058861f
C1835 VDD.t340 VSS 0.013127f
C1836 VDD.n246 VSS 0.059357f
C1837 VDD.t100 VSS 0.05359f
C1838 VDD.t315 VSS 0.05359f
C1839 VDD.t84 VSS 0.070455f
C1840 VDD.n247 VSS 0.081437f
C1841 VDD.t154 VSS 0.082026f
C1842 VDD.t177 VSS 0.068091f
C1843 VDD.t152 VSS 0.068091f
C1844 VDD.t150 VSS 0.081331f
C1845 VDD.n248 VSS 0.032929f
C1846 VDD.t155 VSS 0.0459f
C1847 VDD.n249 VSS 0.088102f
C1848 VDD.n250 VSS 0.034137f
C1849 VDD.n251 VSS 0.081337f
C1850 VDD.t151 VSS 0.0459f
C1851 VDD.n252 VSS 0.065726f
C1852 VDD.n253 VSS 0.055648f
C1853 VDD.n254 VSS 0.089837f
C1854 VDD.t339 VSS 0.08732f
C1855 VDD.n255 VSS 0.086212f
C1856 VDD.n256 VSS 0.039098f
C1857 VDD.t85 VSS 0.038983f
C1858 VDD.n257 VSS 0.085171f
C1859 VDD.t83 VSS 0.038983f
C1860 VDD.n258 VSS 0.085171f
C1861 VDD.n259 VSS 0.039098f
C1862 VDD.n260 VSS 0.086212f
C1863 VDD.t352 VSS 0.070455f
C1864 VDD.t350 VSS 0.05359f
C1865 VDD.t295 VSS 0.05359f
C1866 VDD.t64 VSS 0.05359f
C1867 VDD.t126 VSS 0.05359f
C1868 VDD.t125 VSS 0.05359f
C1869 VDD.t127 VSS 0.05359f
C1870 VDD.t128 VSS 0.05359f
C1871 VDD.t349 VSS 0.05359f
C1872 VDD.t355 VSS 0.05359f
C1873 VDD.t348 VSS 0.05359f
C1874 VDD.t354 VSS 0.05359f
C1875 VDD.t101 VSS 0.05359f
C1876 VDD.t293 VSS 0.05359f
C1877 VDD.t276 VSS 0.05359f
C1878 VDD.t274 VSS 0.071173f
C1879 VDD.n261 VSS 0.083567f
C1880 VDD.n262 VSS 5.68184f
C1881 VDD.t189 VSS 0.078065f
C1882 VDD.n278 VSS 0.050753f
C1883 VDD.n279 VSS 0.172861f
C1884 VDD.t188 VSS 0.061906f
C1885 VDD.n282 VSS 0.084041f
C1886 VDD.t192 VSS 0.044275f
C1887 VDD.n286 VSS 0.084041f
C1888 VDD.t190 VSS 0.044275f
C1889 VDD.n290 VSS 0.084041f
C1890 VDD.t246 VSS 0.044275f
C1891 VDD.t251 VSS 0.077557f
C1892 VDD.n294 VSS 0.1247f
C1893 VDD.n297 VSS 0.125157f
C1894 VDD.t250 VSS 0.072438f
C1895 VDD.n298 VSS 0.084041f
C1896 VDD.n299 VSS 0.048785f
C1897 VDD.t180 VSS 0.014711f
C1898 VDD.t247 VSS 0.014711f
C1899 VDD.n301 VSS 0.051857f
C1900 VDD.n302 VSS 0.028929f
C1901 VDD.n307 VSS 0.048785f
C1902 VDD.t179 VSS 0.044275f
C1903 VDD.n308 VSS 0.084041f
C1904 VDD.n309 VSS 0.048785f
C1905 VDD.t259 VSS 0.014711f
C1906 VDD.t191 VSS 0.014711f
C1907 VDD.n311 VSS 0.051857f
C1908 VDD.n312 VSS 0.028929f
C1909 VDD.n317 VSS 0.048785f
C1910 VDD.t258 VSS 0.044275f
C1911 VDD.n318 VSS 0.084041f
C1912 VDD.n319 VSS 0.048785f
C1913 VDD.t249 VSS 0.014711f
C1914 VDD.t193 VSS 0.014711f
C1915 VDD.n321 VSS 0.051857f
C1916 VDD.n322 VSS 0.028929f
C1917 VDD.n327 VSS 0.048785f
C1918 VDD.t248 VSS 0.044275f
C1919 VDD.n328 VSS 0.084041f
C1920 VDD.n329 VSS 0.048785f
C1921 VDD.n333 VSS 0.789243f
C1922 VDD.n334 VSS 6.555029f
C1923 VDD.n335 VSS 2.19116f
C1924 VDD.n336 VSS 3.1274f
C1925 VDD.n338 VSS 0.083665f
C1926 VDD.n340 VSS 0.051223f
C1927 VDD.n341 VSS 0.078657f
C1928 VDD.n342 VSS 0.093133f
C1929 VDD.n343 VSS 0.093133f
C1930 VDD.n344 VSS 0.083116f
C1931 VDD.n345 VSS 0.052334f
C1932 VDD.n348 VSS 0.02699f
C1933 VDD.t140 VSS 0.026464f
C1934 VDD.n349 VSS 0.091884f
C1935 VDD.n350 VSS 0.35413f
C1936 VDD.n351 VSS 0.35413f
C1937 VDD.n352 VSS 0.03041f
C1938 VDD.n353 VSS 0.032171f
C1939 VDD.t139 VSS 0.237017f
C1940 VDD.n356 VSS 0.032171f
C1941 VDD.n357 VSS 0.018677f
C1942 VDD.n358 VSS 0.035799f
C1943 VDD.n359 VSS 0.060788f
C1944 VDD.n360 VSS 0.040913f
C1945 VDD.n365 VSS 0.021955f
C1946 VDD.n368 VSS 0.419585f
C1947 VDD.t238 VSS 0.188689f
C1948 VDD.t184 VSS 0.13638f
C1949 VDD.t185 VSS 0.13638f
C1950 VDD.t342 VSS 0.13638f
C1951 VDD.t326 VSS 0.13638f
C1952 VDD.t196 VSS 0.13638f
C1953 VDD.t197 VSS 0.13638f
C1954 VDD.t239 VSS 0.13638f
C1955 VDD.t265 VSS 0.13638f
C1956 VDD.t183 VSS 0.102285f
C1957 VDD.n369 VSS 0.06819f
C1958 VDD.t273 VSS 0.102285f
C1959 VDD.t324 VSS 0.13638f
C1960 VDD.t325 VSS 0.13638f
C1961 VDD.t105 VSS 0.13638f
C1962 VDD.t117 VSS 0.13638f
C1963 VDD.t118 VSS 0.13638f
C1964 VDD.t264 VSS 0.13638f
C1965 VDD.t272 VSS 0.13638f
C1966 VDD.t343 VSS 0.13638f
C1967 VDD.t111 VSS 0.188689f
C1968 VDD.n370 VSS 0.419585f
C1969 VDD.n371 VSS 0.013568f
C1970 VDD.n372 VSS 0.051223f
C1971 VDD.n373 VSS 0.133386f
C1972 VDD.n374 VSS 0.115676f
C1973 VDD.n375 VSS 0.051223f
C1974 VDD.n376 VSS 0.093133f
C1975 VDD.n377 VSS 0.093133f
C1976 VDD.n378 VSS 0.088124f
C1977 VDD.n379 VSS 0.094845f
C1978 VDD.n380 VSS 0.419585f
C1979 VDD.t266 VSS 0.188689f
C1980 VDD.t323 VSS 0.13638f
C1981 VDD.t186 VSS 0.13638f
C1982 VDD.t198 VSS 0.13638f
C1983 VDD.t138 VSS 0.13638f
C1984 VDD.t194 VSS 0.13638f
C1985 VDD.t344 VSS 0.13638f
C1986 VDD.t237 VSS 0.13638f
C1987 VDD.t107 VSS 0.13638f
C1988 VDD.t341 VSS 0.102285f
C1989 VDD.n381 VSS 0.06819f
C1990 VDD.t106 VSS 0.102285f
C1991 VDD.t267 VSS 0.13638f
C1992 VDD.t322 VSS 0.13638f
C1993 VDD.t187 VSS 0.13638f
C1994 VDD.t199 VSS 0.13638f
C1995 VDD.t108 VSS 0.13638f
C1996 VDD.t195 VSS 0.13638f
C1997 VDD.t149 VSS 0.13638f
C1998 VDD.t321 VSS 0.13638f
C1999 VDD.t320 VSS 0.188689f
C2000 VDD.n382 VSS 0.419585f
C2001 VDD.n390 VSS 0.040913f
C2002 VDD.n391 VSS 0.229542f
C2003 VDD.n392 VSS 2.6982f
C2004 VDD.t167 VSS 0.101045f
C2005 VDD.n393 VSS 0.107359f
C2006 VDD.t242 VSS 0.101045f
C2007 VDD.n394 VSS 0.112972f
C2008 VDD.n395 VSS 0.066482f
C2009 VDD.n396 VSS 0.742668f
C2010 VDD.n397 VSS 0.869453f
C2011 VDD.n398 VSS 0.011753f
C2012 VDD.t165 VSS 0.101045f
C2013 VDD.n400 VSS 0.067505f
C2014 VDD.t131 VSS 0.140215f
C2015 VDD.n401 VSS 0.140008f
C2016 VDD.n402 VSS 0.011967f
C2017 VDD.n403 VSS 0.099992f
C2018 VDD.n404 VSS 0.553681f
C2019 VDD.n405 VSS 0.011753f
C2020 VDD.t200 VSS 0.101045f
C2021 VDD.n407 VSS 0.067505f
C2022 VDD.t81 VSS 0.140215f
C2023 VDD.n408 VSS 0.140008f
C2024 VDD.n409 VSS 0.011967f
C2025 VDD.n410 VSS 0.099992f
C2026 VDD.n411 VSS 0.553681f
C2027 VDD.n412 VSS 0.011753f
C2028 VDD.t204 VSS 0.101045f
C2029 VDD.n414 VSS 0.067505f
C2030 VDD.t80 VSS 0.140215f
C2031 VDD.n415 VSS 0.140008f
C2032 VDD.n416 VSS 0.011967f
C2033 VDD.n417 VSS 0.099992f
C2034 VDD.n418 VSS 0.553681f
C2035 VDD.n419 VSS 0.011753f
C2036 VDD.t206 VSS 0.101045f
C2037 VDD.n421 VSS 0.067505f
C2038 VDD.t69 VSS 0.140215f
C2039 VDD.n422 VSS 0.140008f
C2040 VDD.n423 VSS 0.011967f
C2041 VDD.n424 VSS 0.099992f
C2042 VDD.n425 VSS 0.553681f
C2043 VDD.n426 VSS 0.011753f
C2044 VDD.t169 VSS 0.101045f
C2045 VDD.n428 VSS 0.067505f
C2046 VDD.t147 VSS 0.140215f
C2047 VDD.n429 VSS 0.140008f
C2048 VDD.n430 VSS 0.011967f
C2049 VDD.n431 VSS 0.099992f
C2050 VDD.n432 VSS 0.553681f
C2051 VDD.n433 VSS 0.011753f
C2052 VDD.t202 VSS 0.101045f
C2053 VDD.n435 VSS 0.067505f
C2054 VDD.t162 VSS 0.140215f
C2055 VDD.n436 VSS 0.140008f
C2056 VDD.n437 VSS 0.011967f
C2057 VDD.n438 VSS 0.099992f
C2058 VDD.n439 VSS 0.457862f
C2059 VDD.n440 VSS 1.1111f
C2060 VDD.n441 VSS 0.022498f
C2061 VDD.t11 VSS 0.075962f
C2062 VDD.t25 VSS 0.117348f
C2063 VDD.t34 VSS 0.117348f
C2064 VDD.t15 VSS 0.117348f
C2065 VDD.t311 VSS 0.124421f
C2066 VDD.t65 VSS 0.076748f
C2067 VDD.t330 VSS 0.094036f
C2068 VDD.t301 VSS 0.053435f
C2069 VDD.t74 VSS 0.077533f
C2070 VDD.t53 VSS 0.091416f
C2071 VDD.t36 VSS 0.072485f
C2072 VDD.n443 VSS 0.240433f
C2073 VDD.n444 VSS 0.033471f
C2074 VDD.n445 VSS 0.036483f
C2075 VDD.n446 VSS 0.037837f
C2076 VDD.n447 VSS 0.040456f
C2077 VDD.n448 VSS 0.042796f
C2078 VDD.n449 VSS 0.040838f
C2079 VDD.n450 VSS 0.040798f
C2080 VDD.n451 VSS 0.035805f
C2081 VDD.n452 VSS 0.033249f
C2082 VDD.n453 VSS 0.040575f
C2083 VDD.n454 VSS 0.037837f
C2084 VDD.n455 VSS 0.026439f
C2085 VDD.n456 VSS 0.032804f
C2086 VDD.n457 VSS 0.037837f
C2087 VDD.n458 VSS 0.034728f
C2088 VDD.n459 VSS 0.024515f
C2089 VDD.n460 VSS 0.037837f
C2090 VDD.n461 VSS 0.040575f
C2091 VDD.n462 VSS 0.021481f
C2092 VDD.n463 VSS 0.035974f
C2093 VDD.n464 VSS 0.123931f
C2094 VDD.t309 VSS 0.0757f
C2095 VDD.t70 VSS 0.071509f
C2096 VDD.t334 VSS 0.099274f
C2097 VDD.t260 VSS 0.09325f
C2098 VDD.t109 VSS 0.100846f
C2099 VDD.t27 VSS 0.069937f
C2100 VDD.t129 VSS 0.09325f
C2101 VDD.t13 VSS 0.117348f
C2102 VDD.t356 VSS 0.053435f
C2103 VDD.t316 VSS 0.117348f
C2104 VDD.t313 VSS 0.11761f
C2105 VDD.t123 VSS 0.09056f
C2106 VDD.n465 VSS 0.027061f
C2107 VDD.n466 VSS 0.255344f
C2108 VDD.n467 VSS 0.399932f
C2109 VDD.n468 VSS 0.031211f
C2110 VDD.n469 VSS 0.203319f
C2111 VDD.t51 VSS 0.079147f
C2112 VDD.t297 VSS 0.117235f
C2113 VDD.t17 VSS 0.117497f
C2114 VDD.t60 VSS 0.06987f
C2115 VDD.t328 VSS 0.100749f
C2116 VDD.t175 VSS 0.09316f
C2117 VDD.t305 VSS 0.099179f
C2118 VDD.t181 VSS 0.07144f
C2119 VDD.t240 VSS 0.09316f
C2120 VDD.t215 VSS 0.117235f
C2121 VDD.t291 VSS 0.053384f
C2122 VDD.t76 VSS 0.08688f
C2123 VDD.n470 VSS 0.112565f
C2124 VDD.t2 VSS 0.075889f
C2125 VDD.t303 VSS 0.08688f
C2126 VDD.n471 VSS 0.123819f
C2127 VDD.t54 VSS 0.084001f
C2128 VDD.t307 VSS 0.061496f
C2129 VDD.t217 VSS 0.106768f
C2130 VDD.t23 VSS 0.062805f
C2131 VDD.t98 VSS 0.053384f
C2132 VDD.t332 VSS 0.053384f
C2133 VDD.t219 VSS 0.062805f
C2134 VDD.t72 VSS 0.068823f
C2135 VDD.n474 VSS 0.081109f
C2136 VDD.t163 VSS 0.062975f
C2137 VDD.n475 VSS 0.082863f
C2138 VDD.n476 VSS 0.259502f
C2139 VDD.n477 VSS 0.042768f
C2140 VDD.n478 VSS 0.017858f
C2141 VDD.n479 VSS 0.033646f
C2142 VDD.n480 VSS 0.037393f
C2143 VDD.n481 VSS 0.034765f
C2144 VDD.n482 VSS 0.035933f
C2145 VDD.n483 VSS 0.023834f
C2146 VDD.n484 VSS 0.05007f
C2147 VDD.n485 VSS 0.040725f
C2148 VDD.n486 VSS 0.033549f
C2149 VDD.n487 VSS 0.021434f
C2150 VDD.n488 VSS 0.040462f
C2151 VDD.n489 VSS 0.037735f
C2152 VDD.n490 VSS 0.026817f
C2153 VDD.n491 VSS 0.032275f
C2154 VDD.n492 VSS 0.037735f
C2155 VDD.n493 VSS 0.035078f
C2156 VDD.n494 VSS 0.024014f
C2157 VDD.n495 VSS 0.037735f
C2158 VDD.n496 VSS 0.040462f
C2159 VDD.n497 VSS 0.033162f
C2160 VDD.n498 VSS 0.025065f
C2161 VDD.n499 VSS 0.0155f
C2162 VDD.n501 VSS 0.013469f
C2163 VDD.n503 VSS 0.031263f
C2164 VDD.n505 VSS 0.634102f
C2165 VDD.n506 VSS 0.031211f
C2166 VDD.t299 VSS 0.090457f
C2167 VDD.t0 VSS 0.122469f
C2168 VDD.t208 VSS 0.162769f
C2169 VDD.t103 VSS 0.166432f
C2170 VDD.t57 VSS 0.150469f
C2171 VDD.t59 VSS 0.081649f
C2172 VDD.n513 VSS 0.100162f
C2173 VDD.t102 VSS 0.058094f
C2174 VDD.t78 VSS 0.095254f
C2175 VDD.t8 VSS 0.134768f
C2176 VDD.t86 VSS 0.152825f
C2177 VDD.t56 VSS 0.115403f
C2178 VDD.t94 VSS 0.105721f
C2179 VDD.t115 VSS 0.155965f
C2180 VDD.t92 VSS 0.18475f
C2181 VDD.n514 VSS 0.10236f
C2182 VDD.t318 VSS 0.307743f
C2183 VDD.n515 VSS 0.095557f
C2184 VDD.n516 VSS 0.099343f
C2185 VDD.n517 VSS 0.030893f
C2186 VDD.n518 VSS 0.051546f
C2187 VDD.n519 VSS 0.073737f
C2188 VDD.n520 VSS 0.107391f
C2189 VDD.n521 VSS 0.149845f
C2190 VDD.n522 VSS 0.105692f
C2191 VDD.n523 VSS 0.065084f
C2192 VDD.n524 VSS 0.04961f
C2193 VDD.n525 VSS 0.022705f
C2194 VDD.n526 VSS 0.0155f
C2195 VDD.n527 VSS 0.011816f
C2196 VDD.n528 VSS 0.255464f
C2197 VDD.n529 VSS 0.038636f
C2198 VDD.n530 VSS 0.463639f
C2199 VDD.n531 VSS 0.031211f
C2200 VDD.t171 VSS 0.090457f
C2201 VDD.t233 VSS 0.189984f
C2202 VDD.t287 VSS 0.063851f
C2203 VDD.t229 VSS 0.086356f
C2204 VDD.t225 VSS 0.053907f
C2205 VDD.t10 VSS 0.039425f
C2206 VDD.t120 VSS 0.058618f
C2207 VDD.t96 VSS 0.109385f
C2208 VDD.t136 VSS 0.068038f
C2209 VDD.t44 VSS 0.053384f
C2210 VDD.t289 VSS 0.058618f
C2211 VDD.t46 VSS 0.068038f
C2212 VDD.t42 VSS 0.103628f
C2213 VDD.t49 VSS 0.058618f
C2214 VDD.t40 VSS 0.037421f
C2215 VDD.n541 VSS 0.130903f
C2216 VDD.t132 VSS 0.019365f
C2217 VDD.t278 VSS 0.039776f
C2218 VDD.t32 VSS 0.062805f
C2219 VDD.t158 VSS 0.056524f
C2220 VDD.t67 VSS 0.053384f
C2221 VDD.t134 VSS 0.078244f
C2222 VDD.t148 VSS 0.063851f
C2223 VDD.t160 VSS 0.069347f
C2224 VDD.t223 VSS 0.068038f
C2225 VDD.t48 VSS 0.046057f
C2226 VDD.t4 VSS 0.058618f
C2227 VDD.t227 VSS 0.064898f
C2228 VDD.t29 VSS 0.053384f
C2229 VDD.t231 VSS 0.070132f
C2230 VDD.t221 VSS 0.084786f
C2231 VDD.t6 VSS 0.053384f
C2232 VDD.t235 VSS 0.095777f
C2233 VDD.n542 VSS 0.070435f
C2234 VDD.n544 VSS 0.090443f
C2235 VDD.n545 VSS 0.015875f
C2236 VDD.n546 VSS 0.05007f
C2237 VDD.n547 VSS 0.037117f
C2238 VDD.n548 VSS 0.040114f
C2239 VDD.n549 VSS 0.028266f
C2240 VDD.n550 VSS 0.037469f
C2241 VDD.n551 VSS 0.068763f
C2242 VDD.n552 VSS 0.044198f
C2243 VDD.n553 VSS 0.039224f
C2244 VDD.n554 VSS 0.045801f
C2245 VDD.n555 VSS 0.044134f
C2246 VDD.n556 VSS 0.039275f
C2247 VDD.n557 VSS 0.031217f
C2248 VDD.n558 VSS 0.04036f
C2249 VDD.n559 VSS 0.029249f
C2250 VDD.n560 VSS 0.031613f
C2251 VDD.n561 VSS 0.022705f
C2252 VDD.n562 VSS 0.011269f
C2253 VDD.n563 VSS 0.011816f
C2254 VDD.n564 VSS 0.255464f
C2255 VDD.n565 VSS 0.038636f
C2256 VDD.n566 VSS 0.621691f
C2257 VDD.n567 VSS 5.61848f
C2258 VDD.n568 VSS 0.455277f
C2259 VDD.n569 VSS 0.067687f
C2260 VDD.n570 VSS 0.016922f
C2261 VDD.n571 VSS 0.016922f
C2262 VDD.n572 VSS 0.016922f
C2263 VDD.n573 VSS 0.067687f
C2264 VDD.n574 VSS 0.067687f
C2265 VDD.n575 VSS 0.067687f
C2266 VDD.n576 VSS 0.016922f
C2267 VDD.n577 VSS 0.016922f
C2268 VDD.n578 VSS 0.016922f
C2269 VDD.n579 VSS 0.067687f
C2270 VDD.n580 VSS 0.067687f
C2271 VDD.n581 VSS 0.065452f
C2272 VDD.n582 VSS 0.016922f
C2273 VDD.n583 VSS 0.016922f
C2274 VDD.n584 VSS 0.036078f
.ends

