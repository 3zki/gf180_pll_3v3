* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt logic_layout F6 DOWN UP GND VDD VCOIN CLK
X0 a_1792_n5184 a_572_n4284.t4 GND.t82 GND.t81 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 a_896_n2729 a_484_n2316.t2 GND.t130 GND.t129 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2 a_1328_n4595 a_896_n4641 VDD.t138 VDD.t137 pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X3 a_3703_68 a_1233_472 a_3519_68 GND.t42 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4 VDD.t163 a_1877_n1888 a_1317_n1888 VDD.t162 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X5 F6.t7 a_1792_n5184 GND.t17 GND.t16 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X6 a_2459_n4595 a_896_n4641 a_1824_n4271 GND.t109 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7 a_1284_n4227 a_484_n4228.t2 GND.t20 GND.t19 nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X8 GND.t80 a_572_n4284.t5 a_484_n3673.t0 GND.t74 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X9 VDD.t45 a_1233_472 a_757_24 VDD.t44 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X10 GND.t112 a_908_n496 a_820_n404 GND.t111 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X11 a_1824_n3709 a_1452_n3665 GND.t146 GND.t113 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X12 GND.t121 a_1356_n496 a_1268_n404 GND.t120 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X13 a_673_n1440 a_224_n1440 VDD.t129 VDD.t128 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X14 a_2704_n3665 a_484_n3673.t2 a_2459_n3297 GND.t45 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X15 a_3703_n1844 a_1233_n1440 a_3519_n1844 GND.t38 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X16 GND.t15 a_1792_n5184 F6.t6 GND.t14 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X17 a_673_472 a_757_24 a_693_68 GND.t50 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X18 a_1452_n3665 a_1332_n3709 a_1284_n3665 GND.t56 nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X19 a_757_n1888.t0 a_3024_n1440 VDD.t23 VDD.t22 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X20 a_693_68 a_224_472 GND.t28 GND.t27 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X21 a_1452_n3665 a_1332_n3709 a_1328_n3297 VDD.t63 pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X22 a_1877_n1888 a_673_n1440 VDD.t96 VDD.t95 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X23 a_1776_n3665 a_896_n3352 a_1452_n3665 GND.t110 nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X24 GND.t54 a_12_n496 a_n76_n404 GND.t53 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X25 a_2576_n1440 a_673_n1440 VDD.t94 VDD.t93 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X26 a_1792_n5184 a_572_n4284.t6 VDD.t88 VDD.t87 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X27 a_1824_n4271 a_1452_n4227 GND.t114 GND.t113 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X28 a_757_24 a_1877_n1888 VDD.t161 VDD.t160 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X29 GND.t13 a_1792_n5184 F6.t5 GND.t12 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X30 VDD.t166 a_1824_n4271 a_1796_n4595 VDD.t165 pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X31 a_2752_n3709 a_2459_n3297 GND.t108 GND.t30 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X32 a_2704_n4227 a_484_n4228.t3 a_2459_n4595 GND.t45 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X33 a_1796_n3297 a_484_n3673.t3 a_1452_n3665 VDD.t48 pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X34 VDD.t17 a_1792_n5184 F6.t15 VDD.t16 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X35 a_896_n3352 a_484_n3673.t4 GND.t131 GND.t46 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X36 F6.t14 a_1792_n5184 VDD.t15 VDD.t14 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X37 a_1452_n4227 a_224_n2800 a_1284_n4227 GND.t56 nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X38 VDD.t43 a_1233_472 a_1877_n1888 VDD.t42 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X39 VDD.t13 a_1792_n5184 F6.t13 VDD.t12 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X40 VDD.t142 a_124_n4756 a_36_n4712 VDD.t141 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X41 a_460_n496 a_372_n404 VDD.t116 VDD.t115 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X42 a_3519_n1844 a_3024_n1440 GND.t24 GND.t23 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X43 GND.t67 a_2752_n3709 a_2704_n3665 GND.t66 nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X44 a_673_472 a_224_472 VDD.t27 VDD.t26 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X45 a_1332_n2408 a_2752_n3709 GND.t65 GND.t64 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X46 a_1824_n3709 a_1452_n3665 VDD.t164 VDD.t20 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X47 a_224_n5184 VCOIN.t0 GND.t126 GND.t125 nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X48 GND.t52 a_2252_n496 a_2164_n404 GND.t51 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X49 a_1776_n4227 a_896_n4641 a_1452_n4227 GND.t110 nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X50 a_1792_n5184 a_572_n4284.t7 GND.t79 GND.t78 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X51 VDD.t110 a_124_n3449 a_36_n3352 VDD.t109 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X52 a_2459_n2683 a_484_n2316.t3 a_1824_n2359 VDD.t123 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X53 a_2752_n4271 a_2459_n4595 GND.t31 GND.t30 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X54 GND.t26 a_1824_n3709 a_1776_n3665 GND.t25 nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X55 GND.t59 a_4044_n2408 a_3956_n2316 GND.t58 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X56 F6.t12 a_1792_n5184 VDD.t11 VDD.t10 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X57 a_2752_n3709 a_2459_n3297 VDD.t119 VDD.t89 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X58 a_1233_n1440 a_673_n1440 VDD.t92 VDD.t91 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X59 F6.t4 a_1792_n5184 GND.t11 GND.t10 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X60 UP.t0 a_757_24 GND.t49 GND.t48 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X61 DOWN.t0 a_757_n1888.t2 GND.t128 GND.t127 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X62 VDD.t135 a_2752_n4271 a_2744_n4595 VDD.t134 pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X63 GND.t119 a_2752_n4271 a_2704_n4227 GND.t66 nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X64 a_3024_472 a_2576_472 VDD.t66 VDD.t65 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X65 a_2744_n4595 a_896_n4641 a_2459_n4595 VDD.t136 pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X66 a_1332_n3709 a_2752_n4271 GND.t118 GND.t64 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X67 VDD.t58 a_757_24 a_673_472 VDD.t57 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X68 a_224_n1440 a_124_n2844 VDD.t33 VDD.t32 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X69 a_124_n3449 a_36_n3352 GND.t94 GND.t93 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X70 a_224_472 CLK.t0 GND.t44 GND.t43 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X71 a_757_24 a_1877_n1888 a_3703_68 GND.t145 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X72 a_2752_n2359 a_2459_n2683 VDD.t90 VDD.t89 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X73 GND.t147 a_1824_n4271 a_1776_n4227 GND.t25 nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X74 a_2576_472 a_673_472 GND.t99 GND.t98 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X75 a_1317_n1888 a_1233_n1440 VDD.t39 VDD.t38 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X76 a_1328_n2683 a_896_n2729 VDD.t146 VDD.t121 pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X77 VDD.t154 a_224_n5184 a_572_n4284.t1 VDD.t153 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X78 a_896_n4641 a_484_n4228.t4 VDD.t50 VDD.t49 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X79 a_896_n3352 a_484_n3673.t5 VDD.t145 VDD.t124 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X80 a_757_n1888.t0 a_1877_n1888 VDD.t159 VDD.t158 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X81 a_2459_n2683 a_896_n2729 a_1824_n2359 GND.t133 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X82 a_1284_n2315 a_484_n2316.t4 GND.t124 GND.t123 nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X83 a_1877_n1888 a_1233_472 a_3473_n404 GND.t41 nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X84 VDD.t9 a_1792_n5184 F6.t11 VDD.t8 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X85 a_693_n1844 a_224_n1440 GND.t116 GND.t115 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X86 a_1452_n4227 a_224_n2800 a_1328_n4595 VDD.t155 pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X87 a_124_n4756 a_36_n4712 GND.t117 GND.t93 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X88 GND.t77 a_572_n4284.t8 a_1792_n5184 GND.t76 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X89 GND.t75 a_572_n4284.t9 a_484_n4228.t0 GND.t74 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X90 a_3519_68 a_3024_472 GND.t1 GND.t0 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X91 a_3024_n1440 a_2576_n1440 VDD.t107 VDD.t106 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X92 a_1317_24 a_1233_472 VDD.t41 VDD.t40 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X93 a_896_n2729 a_484_n2316.t5 VDD.t125 VDD.t124 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X94 a_2459_n3297 a_484_n3673.t6 a_1824_n3709 VDD.t123 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X95 GND.t107 a_460_n496 a_372_n404 GND.t106 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X96 a_1317_24 a_1877_n1888 a_1813_68 GND.t144 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X97 a_572_n4284.t1 a_224_n5184 VDD.t152 VDD.t151 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X98 a_1233_472 a_673_472 VDD.t105 VDD.t104 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X99 a_1813_68 a_1233_472 GND.t40 GND.t39 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X100 a_1796_n4595 a_484_n4228.t5 a_1452_n4227 VDD.t99 pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X101 a_1824_n2359 a_1452_n2315 GND.t22 GND.t21 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X102 a_224_n2800 a_124_n2844 VDD.t31 VDD.t30 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X103 F6.t10 a_1792_n5184 VDD.t7 VDD.t6 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X104 a_1804_n496 a_1716_n404 VDD.t52 VDD.t51 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X105 VDD.t64 a_1824_n2359 a_1796_n2683 VDD.t24 pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X106 a_224_n5184 VCOIN.t1 VDD.t140 VDD.t139 pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X107 a_673_n1440 a_757_n1888.t3 a_693_n1844 GND.t102 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X108 a_2704_n2315 a_484_n2316.t6 a_2459_n2683 GND.t29 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X109 a_1452_n2315 a_1332_n2408 a_1284_n2315 GND.t57 nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X110 VDD.t150 a_224_n5184 a_572_n4284.t0 VDD.t149 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X111 a_1332_n3709 a_2752_n4271 VDD.t133 VDD.t132 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X112 a_1824_n4271 a_1452_n4227 VDD.t127 VDD.t126 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X113 a_2576_n1440 a_673_n1440 GND.t90 GND.t89 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X114 a_896_n4641 a_484_n4228.t6 GND.t47 GND.t46 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X115 VDD.t157 a_1877_n1888 a_1317_24 VDD.t156 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X116 a_1776_n2315 a_896_n2729 a_1452_n2315 GND.t132 nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X117 a_1332_n2408 a_2752_n3709 VDD.t71 VDD.t70 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X118 a_1328_n3297 a_896_n3352 VDD.t122 VDD.t121 pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X119 VDD.t114 a_1317_24 a_1233_472 VDD.t113 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X120 a_3473_n404 a_673_472 a_3269_n404 GND.t97 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X121 a_2752_n2359 a_2459_n2683 GND.t84 GND.t83 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X122 a_4044_n4320 a_3956_n4228 VDD.t112 VDD.t111 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X123 F6.t3 a_1792_n5184 GND.t9 GND.t8 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X124 VDD.t98 a_757_n1888.t4 a_673_n1440 VDD.t97 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X125 a_757_n1888.t1 a_1877_n1888 a_3703_n1844 GND.t143 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X126 VDD.t144 VCOIN.t2 a_224_n5184 VDD.t143 pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X127 VDD.t47 a_4044_n3449 a_3956_n3352 VDD.t46 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X128 a_1253_n1844 a_673_n1440 GND.t88 GND.t87 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X129 GND.t141 a_224_n5184 a_572_n4284.t2 GND.t140 nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X130 a_572_n4284.t0 a_224_n5184 VDD.t148 VDD.t147 pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X131 a_1877_n1888 a_673_472 VDD.t103 VDD.t102 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X132 GND.t71 a_2752_n2359 a_2704_n2315 GND.t70 nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X133 VDD.t75 a_2752_n2359 a_2744_n2683 VDD.t68 pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X134 a_757_24 a_3024_472 VDD.t1 VDD.t0 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X135 a_124_n2844 a_2752_n2359 GND.t69 GND.t68 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X136 a_2744_n2683 a_896_n2729 a_2459_n2683 VDD.t120 pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X137 a_1233_472 a_1317_24 a_1253_68 GND.t105 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X138 a_1253_68 a_673_472 GND.t96 GND.t95 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X139 a_908_n496 a_820_n404 VDD.t60 VDD.t59 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X140 a_1356_n496 a_1268_n404 VDD.t54 VDD.t53 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X141 GND.t61 a_1824_n2359 a_1776_n2315 GND.t60 nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X142 F6.t2 a_1792_n5184 GND.t7 GND.t6 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X143 a_3075_n404 a_673_n1440 GND.t86 GND.t85 nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X144 a_1813_n1844 a_1233_n1440 GND.t37 GND.t36 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X145 a_4044_n3449 a_3956_n3352 GND.t92 GND.t91 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X146 VDD.t86 a_572_n4284.t10 a_484_n3673.t1 VDD.t80 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X147 VDD.t83 a_572_n4284.t11 a_1792_n5184 VDD.t82 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X148 VDD.t85 a_572_n4284.t12 a_484_n4228.t1 VDD.t84 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X149 VDD.t37 a_1233_n1440 a_757_n1888.t0 VDD.t36 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X150 a_1233_n1440 a_1317_n1888 a_1253_n1844 GND.t18 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X151 a_224_n1440 a_124_n2844 GND.t34 GND.t32 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X152 VDD.t25 a_1824_n3709 a_1796_n3297 VDD.t24 pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X153 a_3024_472 a_2576_472 GND.t63 GND.t62 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X154 GND.t5 a_1792_n5184 F6.t1 GND.t4 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X155 a_572_n4284.t2 a_224_n5184 GND.t139 GND.t138 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X156 F6.t9 a_1792_n5184 VDD.t5 VDD.t4 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X157 UP.t1 a_757_24 VDD.t56 VDD.t55 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X158 a_12_n496 a_n76_n404 VDD.t62 VDD.t61 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X159 a_224_n2800 a_124_n2844 GND.t33 GND.t32 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X160 a_1452_n2315 a_1332_n2408 a_1328_n2683 VDD.t63 pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X161 GND.t104 a_1804_n496 a_1716_n404 GND.t103 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X162 DOWN.t1 a_757_n1888.t5 VDD.t73 VDD.t72 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X163 GND.t73 a_572_n4284.t13 a_484_n2316.t0 GND.t72 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X164 a_2459_n4595 a_484_n4228.t7 a_1824_n4271 VDD.t108 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X165 GND.t137 a_224_n5184 a_572_n4284.t3 GND.t136 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X166 a_224_472 CLK.t1 VDD.t131 VDD.t130 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X167 VDD.t81 a_572_n4284.t14 a_484_n2316.t1 VDD.t80 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X168 VDD.t79 a_572_n4284.t15 a_1792_n5184 VDD.t78 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X169 a_1317_n1888 a_1877_n1888 a_1813_n1844 GND.t142 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X170 GND.t122 a_4044_n4320 a_3956_n4228 GND.t91 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X171 a_3269_n404 a_1233_n1440 a_3075_n404 GND.t35 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X172 GND.t3 a_1792_n5184 F6.t0 GND.t2 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X173 a_1792_n5184 a_572_n4284.t16 VDD.t77 VDD.t76 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X174 a_2576_472 a_673_472 VDD.t101 VDD.t100 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X175 a_124_n2844 a_2752_n2359 VDD.t74 VDD.t70 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X176 VDD.t19 a_1317_n1888 a_1233_n1440 VDD.t18 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X177 a_1796_n2683 a_484_n2316.t7 a_1452_n2315 VDD.t48 pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X178 VDD.t3 a_1792_n5184 F6.t8 VDD.t2 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X179 a_2459_n3297 a_896_n3352 a_1824_n3709 GND.t109 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X180 a_2252_n496 a_2164_n404 VDD.t118 VDD.t117 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X181 a_1284_n3665 a_484_n3673.t7 GND.t55 GND.t19 nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X182 VDD.t35 a_1233_n1440 a_1877_n1888 VDD.t34 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X183 a_3024_n1440 a_2576_n1440 GND.t101 GND.t100 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X184 VDD.t69 a_2752_n3709 a_2744_n3297 VDD.t68 pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X185 a_1824_n2359 a_1452_n2315 VDD.t21 VDD.t20 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X186 a_2752_n4271 a_2459_n4595 VDD.t29 VDD.t28 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X187 a_2744_n3297 a_896_n3352 a_2459_n3297 VDD.t120 pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X188 a_4044_n2408 a_3956_n2316 VDD.t67 VDD.t46 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X189 a_572_n4284.t3 a_224_n5184 GND.t135 GND.t134 nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
R0 a_572_n4284.n2 a_572_n4284.t11 31.6987
R1 a_572_n4284.n3 a_572_n4284.t16 18.6885
R2 a_572_n4284.n0 a_572_n4284.t15 18.6885
R3 a_572_n4284.n2 a_572_n4284.t6 18.6885
R4 a_572_n4284.n5 a_572_n4284.t5 13.907
R5 a_572_n4284.n4 a_572_n4284.t13 13.8462
R6 a_572_n4284.n6 a_572_n4284.t9 13.8462
R7 a_572_n4284.n4 a_572_n4284.t14 12.1185
R8 a_572_n4284.n6 a_572_n4284.t12 12.1185
R9 a_572_n4284.n5 a_572_n4284.t10 12.0455
R10 a_572_n4284.n3 a_572_n4284.t4 11.1938
R11 a_572_n4284.n0 a_572_n4284.t8 11.1938
R12 a_572_n4284.n2 a_572_n4284.t7 11.1938
R13 a_572_n4284.n1 a_572_n4284.n4 10.6383
R14 a_572_n4284.n0 a_572_n4284.n3 10.5449
R15 a_572_n4284.n1 a_572_n4284.n6 10.2813
R16 a_572_n4284.n1 a_572_n4284.n5 10.2813
R17 a_572_n4284.n0 a_572_n4284.n1 8.87498
R18 a_572_n4284.n0 a_572_n4284.t3 7.33746
R19 a_572_n4284.n0 a_572_n4284.n2 6.48939
R20 a_572_n4284.n0 a_572_n4284.t2 6.46093
R21 a_572_n4284.t0 a_572_n4284.n0 6.01368
R22 a_572_n4284.n0 a_572_n4284.t1 5.4118
R23 GND.n83 GND.n82 19865.5
R24 GND.n62 GND.n6 18793.3
R25 GND.n82 GND.n62 17721.1
R26 GND.t78 GND.t6 3591.32
R27 GND.t125 GND.t134 3591.32
R28 GND.t140 GND.t81 3057.08
R29 GND.n83 GND.t125 2226.03
R30 GND.t72 GND.t32 1662.1
R31 GND.t10 GND.t14 1662.1
R32 GND.t12 GND.t10 1662.1
R33 GND.t16 GND.t12 1662.1
R34 GND.t4 GND.t16 1662.1
R35 GND.t8 GND.t4 1662.1
R36 GND.t2 GND.t8 1662.1
R37 GND.t6 GND.t2 1662.1
R38 GND.t76 GND.t78 1662.1
R39 GND.t81 GND.t76 1662.1
R40 GND.t138 GND.t140 1662.1
R41 GND.t136 GND.t138 1662.1
R42 GND.t134 GND.t136 1662.1
R43 GND.t74 GND.t93 1513.7
R44 GND.t64 GND.t30 1439.5
R45 GND.t23 GND.t83 1406.11
R46 GND.t106 GND.t43 1394.98
R47 GND.t19 GND.t46 1365.3
R48 GND.n81 GND.t93 1261.42
R49 GND.t87 GND.t129 1250.29
R50 GND.n69 GND.t64 1246.58
R51 GND.n72 GND.t91 1231.74
R52 GND.t132 GND.t57 1202.05
R53 GND.t110 GND.t56 1202.05
R54 GND.t113 GND.t25 1157.53
R55 GND.n14 GND.t62 1113.01
R56 GND.n61 GND.t32 1113.01
R57 GND.n15 GND.t144 1109.3
R58 GND.t39 GND.t120 1101.88
R59 GND.t143 GND.t58 1101.88
R60 GND.n62 GND.n61 1072.2
R61 GND.n82 GND.n81 1072.2
R62 GND.t30 GND.t66 994.293
R63 GND.t21 GND.t142 960.903
R64 GND.t53 GND.n6 845.89
R65 GND.n34 GND.n33 831.051
R66 GND.t45 GND.t109 831.051
R67 GND.t109 GND.t113 831.051
R68 GND.t46 GND.t74 831.051
R69 GND.t42 GND.t145 756.85
R70 GND.t35 GND.t97 756.85
R71 GND.t85 GND.t35 719.75
R72 GND.t111 GND.t50 708.62
R73 GND.t95 GND.t111 686.359
R74 GND.t51 GND.t98 682.649
R75 GND.t105 GND.t95 682.649
R76 GND.t50 GND.t27 682.649
R77 GND.t133 GND.n9 682.649
R78 GND.t102 GND.t115 682.649
R79 GND.t38 GND.t68 649.259
R80 GND.t100 GND.t70 638.129
R81 GND.n46 GND.t38 626.999
R82 GND.t70 GND.t29 623.288
R83 GND.t66 GND.t45 623.288
R84 GND.t25 GND.t110 623.288
R85 GND.t56 GND.t19 623.288
R86 GND.t18 GND.t123 567.638
R87 GND.t103 GND.t39 560.217
R88 GND.t48 GND.n12 554.422
R89 GND.t0 GND.t41 549.087
R90 GND.t98 GND.n14 549.087
R91 GND.t60 GND.t36 486.017
R92 GND.n15 GND.t51 430.365
R93 GND.t89 GND.t133 430.365
R94 GND.t29 GND.t89 400.685
R95 GND.t83 GND.t100 356.164
R96 GND.t120 GND.t105 293.094
R97 GND.n34 GND.t48 281.964
R98 GND.t27 GND.t106 270.834
R99 GND.t43 GND.t53 267.123
R100 GND.t58 GND.t127 267.123
R101 GND.n33 GND.t145 255.994
R102 GND.t142 GND.t60 196.632
R103 GND.t97 GND.t0 170.662
R104 GND.n9 GND.t21 148.403
R105 GND.t129 GND.t102 144.692
R106 GND.t36 GND.t132 137.273
R107 GND.t41 GND.t42 133.562
R108 GND.n46 GND.t143 129.852
R109 GND.t144 GND.t103 122.433
R110 GND.t62 GND.t85 115.011
R111 GND.t123 GND.t87 115.011
R112 GND.t57 GND.t18 55.6512
R113 GND.t68 GND.t23 33.3909
R114 GND.n72 GND.n69 29.6809
R115 GND.n54 GND.n8 12.033
R116 GND.n77 GND.n66 12.033
R117 GND.n77 GND.n65 12.033
R118 GND.n56 GND.t124 11.0292
R119 GND.n78 GND.t20 11.0292
R120 GND.n78 GND.t55 11.0292
R121 GND.n88 GND.t82 10.5091
R122 GND.n94 GND.t15 10.3593
R123 GND.n90 GND.t7 10.2792
R124 GND.n87 GND.t141 10.0514
R125 GND.n85 GND.t135 10.0514
R126 GND.n35 GND.t49 9.93604
R127 GND.n29 GND.t63 9.93604
R128 GND.n26 GND.t99 9.93604
R129 GND.n16 GND.t44 9.93604
R130 GND.n11 GND.t128 9.93604
R131 GND.n51 GND.t101 9.93604
R132 GND.n52 GND.t90 9.93604
R133 GND.n60 GND.t33 9.93604
R134 GND.n60 GND.t34 9.93604
R135 GND.n84 GND.t126 9.15882
R136 GND.n70 GND.t122 8.53771
R137 GND.n42 GND.t59 8.51229
R138 GND.n17 GND.t54 8.51132
R139 GND.n19 GND.t107 8.51132
R140 GND.n21 GND.t112 8.51132
R141 GND.n22 GND.t121 8.51132
R142 GND.n24 GND.t104 8.51132
R143 GND.n27 GND.t52 8.51132
R144 GND.n71 GND.t92 8.51132
R145 GND.n80 GND.t117 8.51132
R146 GND.n80 GND.t94 8.51132
R147 GND.n30 GND.t86 8.48197
R148 GND.n48 GND.t69 8.46241
R149 GND.n75 GND.t118 8.46241
R150 GND.n75 GND.t65 8.46241
R151 GND.n31 GND.t1 8.4135
R152 GND.n23 GND.t40 8.4135
R153 GND.n20 GND.t96 8.4135
R154 GND.n18 GND.t28 8.4135
R155 GND.n49 GND.t24 8.4135
R156 GND.n55 GND.t37 8.4135
R157 GND.n57 GND.t88 8.4135
R158 GND.n59 GND.t116 8.4135
R159 GND.n8 GND.t22 8.4005
R160 GND.n8 GND.t61 8.4005
R161 GND.n66 GND.t114 8.4005
R162 GND.n66 GND.t147 8.4005
R163 GND.n65 GND.t146 8.4005
R164 GND.n65 GND.t26 8.4005
R165 GND.n10 GND.t71 8.0855
R166 GND.n68 GND.t119 8.0855
R167 GND.n67 GND.t67 8.0855
R168 GND.n50 GND.n10 6.54898
R169 GND.n76 GND.n67 6.54898
R170 GND.n76 GND.n68 6.54898
R171 GND.n58 GND.n7 6.46859
R172 GND.n79 GND.n63 6.46859
R173 GND.n79 GND.n64 6.46859
R174 GND.n89 GND.n4 6.46462
R175 GND.n93 GND.n1 6.45138
R176 GND.n92 GND.n2 6.45138
R177 GND.n91 GND.n3 6.45138
R178 GND.n86 GND.n5 6.45138
R179 GND.n84 GND.n83 5.46326
R180 GND.n16 GND.n6 5.38021
R181 GND.n28 GND.n14 5.32359
R182 GND.n33 GND.n32 5.32359
R183 GND.n36 GND.n34 5.32359
R184 GND.n47 GND.n46 5.32359
R185 GND.n73 GND.n72 5.32359
R186 GND.n25 GND.n15 5.32226
R187 GND.n53 GND.n9 5.32226
R188 GND.n74 GND.n69 5.32226
R189 GND.n10 GND.t84 4.0955
R190 GND.n68 GND.t31 4.0955
R191 GND.n67 GND.t108 4.0955
R192 GND.n4 GND.t79 4.04494
R193 GND.n4 GND.t77 4.04494
R194 GND.n7 GND.t130 4.04494
R195 GND.n7 GND.t73 4.04494
R196 GND.n64 GND.t47 4.04494
R197 GND.n64 GND.t75 4.04494
R198 GND.n63 GND.t131 4.04494
R199 GND.n63 GND.t80 4.04494
R200 GND.n1 GND.t11 3.8098
R201 GND.n1 GND.t13 3.8098
R202 GND.n2 GND.t17 3.8098
R203 GND.n2 GND.t5 3.8098
R204 GND.n3 GND.t9 3.8098
R205 GND.n3 GND.t3 3.8098
R206 GND.t115 GND.t72 3.71055
R207 GND.n5 GND.t139 3.6005
R208 GND.n5 GND.t137 3.6005
R209 GND.n61 GND.n60 2.72066
R210 GND.n81 GND.n80 2.72066
R211 GND.n38 GND.n13 2.28317
R212 GND.n45 GND.n44 2.28317
R213 GND.n38 GND.n37 2.2505
R214 GND.n44 GND.n43 2.2505
R215 GND.n95 GND.n94 2.23903
R216 GND.n42 GND.n41 1.15798
R217 GND.n39 GND.n12 1.14765
R218 GND.n70 GND.n0 1.12597
R219 GND.n40 GND.n39 0.9215
R220 GND.n41 GND.n40 0.563
R221 GND.n90 GND.n89 0.3635
R222 GND.n85 GND.n84 0.3635
R223 GND.n40 GND.n0 0.359
R224 GND.n95 GND.n0 0.342875
R225 GND.n93 GND.n92 0.3365
R226 GND.n92 GND.n91 0.3365
R227 GND.n91 GND.n90 0.3365
R228 GND.n89 GND.n88 0.3365
R229 GND.n87 GND.n86 0.3365
R230 GND.n86 GND.n85 0.3365
R231 GND.n77 GND.n76 0.286527
R232 GND.n78 GND.n77 0.286527
R233 GND.n94 GND.n93 0.235423
R234 GND.n80 GND.n79 0.207623
R235 GND.n32 GND.n31 0.175877
R236 GND.n56 GND.n55 0.163548
R237 GND.n88 GND.n87 0.1415
R238 GND.n48 GND.n47 0.141048
R239 GND.n60 GND.n59 0.13889
R240 GND.n22 GND.n21 0.138582
R241 GND.n52 GND.n51 0.138582
R242 GND.n75 GND.n74 0.138582
R243 GND.n31 GND.n30 0.137349
R244 GND.n24 GND.n23 0.128411
R245 GND.n55 GND.n54 0.123479
R246 GND.n76 GND.n75 0.120089
R247 GND.n50 GND.n49 0.117315
R248 GND.n20 GND.n19 0.114233
R249 GND.n79 GND.n78 0.113925
R250 GND.n58 GND.n57 0.10437
R251 GND.n47 GND.n45 0.083411
R252 GND.n18 GND.n17 0.0797123
R253 GND.n71 GND.n70 0.0704815
R254 GND.n59 GND.n58 0.0692329
R255 GND.n54 GND.n53 0.060911
R256 GND.n17 GND.n16 0.0596781
R257 GND.n19 GND.n18 0.0593699
R258 GND.n29 GND.n28 0.0584452
R259 GND.n26 GND.n25 0.0584452
R260 GND.n53 GND.n52 0.0584452
R261 GND.n28 GND.n27 0.0559795
R262 GND.n25 GND.n24 0.0559795
R263 GND.n73 GND.n71 0.0559795
R264 GND.n32 GND.n13 0.0513562
R265 GND.n37 GND.n12 0.0444564
R266 GND.n43 GND.n42 0.0341269
R267 GND.n51 GND.n50 0.030089
R268 GND.n43 GND.n11 0.0260822
R269 GND.n27 GND.n26 0.0251575
R270 GND.n21 GND.n20 0.0248493
R271 GND.n39 GND.n38 0.0168356
R272 GND.n44 GND.n41 0.0168356
R273 GND.n37 GND.n36 0.0149863
R274 GND.n36 GND.n35 0.0115959
R275 GND GND.n95 0.011375
R276 GND.n23 GND.n22 0.0106712
R277 GND.n30 GND.n29 0.0100548
R278 GND.n57 GND.n56 0.0100548
R279 GND.n35 GND.n13 0.00758904
R280 GND.n45 GND.n11 0.00758904
R281 GND.n49 GND.n48 0.00327397
R282 GND.n74 GND.n73 0.00296575
R283 a_484_n2316.n2 a_484_n2316.t3 121.874
R284 a_484_n2316.t3 a_484_n2316.t6 61.5152
R285 a_484_n2316.n0 a_484_n2316.t4 52.378
R286 a_484_n2316.n0 a_484_n2316.t5 17.7882
R287 a_484_n2316.n1 a_484_n2316.t0 11.1158
R288 a_484_n2316.n1 a_484_n2316.n2 9.95623
R289 a_484_n2316.n1 a_484_n2316.n0 8.37615
R290 a_484_n2316.t1 a_484_n2316.n1 8.02846
R291 a_484_n2316.n0 a_484_n2316.t2 7.3005
R292 a_484_n2316.n2 a_484_n2316.t7 6.7165
R293 VDD.t65 VDD.t0 916.989
R294 VDD.t130 VDD.t26 866.795
R295 VDD.t100 VDD.t65 864.865
R296 VDD.t113 VDD.t40 687.26
R297 VDD.t57 VDD.t104 687.26
R298 VDD.t160 VDD.t55 673.745
R299 VDD.n115 VDD.t130 564.235
R300 VDD.n114 VDD.t100 559.846
R301 VDD.t156 VDD.n114 557.915
R302 VDD.t121 VDD.t124 416.988
R303 VDD.t80 VDD.t109 403.476
R304 VDD.t44 VDD.t160 393.822
R305 VDD.t0 VDD.t44 393.822
R306 VDD.t40 VDD.t156 393.822
R307 VDD.t104 VDD.t113 393.822
R308 VDD.t26 VDD.t57 393.822
R309 VDD.t115 VDD.t32 372.587
R310 VDD.n43 VDD.t70 345.56
R311 VDD.t70 VDD.t89 335.908
R312 VDD.n44 VDD.t46 320.464
R313 VDD.t123 VDD.t20 288.611
R314 VDD.n33 VDD.t139 282.116
R315 VDD.n57 VDD.t30 282.116
R316 VDD.t106 VDD.n63 279.923
R317 VDD.n62 VDD.t162 278.959
R318 VDD.t38 VDD.t53 277.027
R319 VDD.t120 VDD.t123 275.098
R320 VDD.t89 VDD.t68 239.382
R321 VDD.t16 VDD.t14 235.522
R322 VDD.t84 VDD.t143 235.522
R323 VDD.n11 VDD.t6 233.591
R324 VDD.t10 VDD.t82 231.661
R325 VDD.t61 VDD.n61 224.436
R326 VDD.n67 VDD.n66 217.452
R327 VDD.t151 VDD.t149 216.216
R328 VDD.t108 VDD.t87 211.391
R329 VDD.t20 VDD.t24 208.494
R330 VDD.t158 VDD.t36 196.911
R331 VDD.t102 VDD.t34 196.911
R332 VDD.t34 VDD.t95 196.911
R333 VDD.t18 VDD.t91 196.911
R334 VDD.t97 VDD.t128 196.911
R335 VDD.t124 VDD.t80 196.911
R336 VDD.t12 VDD.t4 196.911
R337 VDD.t49 VDD.t147 181.468
R338 VDD.t59 VDD.t97 174.71
R339 VDD.t28 VDD.t2 173.745
R340 VDD.t91 VDD.t59 168.919
R341 VDD.t93 VDD.t117 167.954
R342 VDD.t143 VDD.t141 167.954
R343 VDD.t137 VDD.t151 166.024
R344 VDD.t42 VDD.t22 162.162
R345 VDD.t51 VDD.t38 155.405
R346 VDD.n63 VDD.t93 152.511
R347 VDD.t68 VDD.t120 150.579
R348 VDD.t134 VDD.t136 150.579
R349 VDD.t24 VDD.t48 142.857
R350 VDD.t165 VDD.t99 142.857
R351 VDD.n42 VDD.t121 138.031
R352 VDD.t4 VDD.t111 121.623
R353 VDD.t6 VDD.t132 119.692
R354 VDD.t126 VDD.t78 119.692
R355 VDD.t111 VDD.t8 113.9
R356 VDD.t117 VDD.n62 111.969
R357 VDD.t78 VDD.t165 88.8036
R358 VDD.n10 VDD.t153 87.8383
R359 VDD.t132 VDD.t16 77.2206
R360 VDD.t87 VDD.t126 77.2206
R361 VDD.t48 VDD.n42 71.4291
R362 VDD.t76 VDD.n10 67.5681
R363 VDD.t53 VDD.t18 66.6028
R364 VDD.t2 VDD.t134 65.6376
R365 VDD.t128 VDD.t115 60.8113
R366 VDD.t32 VDD.t61 59.8461
R367 VDD.n66 VDD.t158 56.9503
R368 VDD.t153 VDD.t137 50.1936
R369 VDD.t109 VDD.t30 48.263
R370 VDD.t141 VDD.t139 48.263
R371 VDD.n67 VDD.t72 44.4358
R372 VDD.t162 VDD.t51 41.5063
R373 VDD.t36 VDD.t42 34.7495
R374 VDD.t22 VDD.t102 34.7495
R375 VDD.t149 VDD.t49 34.7495
R376 VDD.t95 VDD.t106 29.9233
R377 VDD.t82 VDD.t108 24.1318
R378 VDD.t14 VDD.t28 23.1665
R379 VDD.n51 VDD.t122 21.6375
R380 VDD.n51 VDD.t146 21.6375
R381 VDD.n25 VDD.t138 21.6375
R382 VDD.t136 VDD.t10 19.3055
R383 VDD.n10 VDD.t155 16.2012
R384 VDD.n42 VDD.t63 15.981
R385 VDD.t147 VDD.t84 15.4445
R386 VDD.n44 VDD.n43 7.72251
R387 VDD.n31 VDD.t140 7.51784
R388 VDD.n23 VDD.t77 7.5061
R389 VDD.n71 VDD.t43 7.46
R390 VDD.n74 VDD.t96 7.46
R391 VDD.n41 VDD.t69 7.40883
R392 VDD.n40 VDD.t75 7.40883
R393 VDD.n7 VDD.t135 7.40883
R394 VDD.n39 VDD.t25 6.22272
R395 VDD.n38 VDD.t64 6.22272
R396 VDD.n4 VDD.t166 6.22272
R397 VDD.n49 VDD.n40 5.49789
R398 VDD.n49 VDD.n41 5.49789
R399 VDD.n19 VDD.n7 5.49789
R400 VDD.n50 VDD.n38 5.41359
R401 VDD.n50 VDD.n39 5.41359
R402 VDD.n22 VDD.n4 5.41359
R403 VDD.n26 VDD.n3 5.35702
R404 VDD.n21 VDD.n5 5.35702
R405 VDD.n18 VDD.n8 5.35702
R406 VDD.n16 VDD.n9 5.35702
R407 VDD.n14 VDD.n12 5.35702
R408 VDD.n52 VDD.n36 5.35271
R409 VDD.n52 VDD.n37 5.35271
R410 VDD.n27 VDD.n2 5.35271
R411 VDD.n28 VDD.n1 5.31398
R412 VDD.n73 VDD.n64 5.30615
R413 VDD.n101 VDD.n100 5.29976
R414 VDD.n70 VDD.n65 5.29976
R415 VDD.n20 VDD.n6 5.28659
R416 VDD.n39 VDD.t164 5.05606
R417 VDD.n38 VDD.t21 5.05606
R418 VDD.n4 VDD.t127 5.05606
R419 VDD.n102 VDD.t1 4.70061
R420 VDD.n72 VDD.t23 4.70061
R421 VDD.n101 VDD.t56 4.62601
R422 VDD.n106 VDD.n98 4.58
R423 VDD.n99 VDD.n98 4.5005
R424 VDD.n107 VDD.t27 4.46351
R425 VDD.n108 VDD.t58 4.46351
R426 VDD.n109 VDD.t105 4.46351
R427 VDD.n110 VDD.t114 4.46351
R428 VDD.n111 VDD.t41 4.46351
R429 VDD.n112 VDD.t157 4.46351
R430 VDD.n88 VDD.t129 4.46351
R431 VDD.n86 VDD.t98 4.46351
R432 VDD.n85 VDD.t92 4.46351
R433 VDD.n83 VDD.t19 4.46351
R434 VDD.n82 VDD.t39 4.46351
R435 VDD.n80 VDD.t163 4.46351
R436 VDD.n45 VDD.t47 4.45405
R437 VDD.n13 VDD.t9 4.385
R438 VDD.n105 VDD.t131 4.36426
R439 VDD.n104 VDD.t101 4.36426
R440 VDD.n103 VDD.t66 4.36426
R441 VDD.n91 VDD.t33 4.36426
R442 VDD.n77 VDD.t94 4.36426
R443 VDD.n75 VDD.t107 4.36426
R444 VDD.n68 VDD.t73 4.36426
R445 VDD.n55 VDD.t31 4.36426
R446 VDD.n79 VDD.t118 4.36035
R447 VDD.n81 VDD.t52 4.36035
R448 VDD.n84 VDD.t54 4.36035
R449 VDD.n87 VDD.t60 4.36035
R450 VDD.n89 VDD.t116 4.36035
R451 VDD.n93 VDD.t62 4.36035
R452 VDD.n45 VDD.t67 4.36035
R453 VDD.n53 VDD.t110 4.36035
R454 VDD.n13 VDD.t112 4.36035
R455 VDD.n29 VDD.t142 4.36035
R456 VDD.n114 VDD.n113 4.35926
R457 VDD.n78 VDD.n62 4.35926
R458 VDD.n47 VDD.n43 4.35926
R459 VDD.n69 VDD.n66 4.35925
R460 VDD.n76 VDD.n63 4.35925
R461 VDD.n46 VDD.n44 4.35925
R462 VDD.n15 VDD.n11 4.35925
R463 VDD.n48 VDD.t71 4.29774
R464 VDD.n48 VDD.t74 4.29774
R465 VDD.n17 VDD.t133 4.29774
R466 VDD.n24 VDD.t154 4.28209
R467 VDD.n1 VDD.t148 3.91054
R468 VDD.t99 VDD.t76 3.8615
R469 VDD.n6 VDD.t83 3.7566
R470 VDD.n68 VDD.n67 3.05229
R471 VDD.n116 VDD.n115 2.3007
R472 VDD.n95 VDD.n61 2.29149
R473 VDD.n90 VDD.n60 2.28317
R474 VDD.n54 VDD.n35 2.28317
R475 VDD.n30 VDD.n0 2.28317
R476 VDD.n41 VDD.t119 2.2755
R477 VDD.n40 VDD.t90 2.2755
R478 VDD.n7 VDD.t29 2.2755
R479 VDD.n95 VDD.n94 2.2505
R480 VDD.n92 VDD.n60 2.2505
R481 VDD.n56 VDD.n35 2.2505
R482 VDD.n32 VDD.n0 2.2505
R483 VDD.n1 VDD.t144 2.22001
R484 VDD.n5 VDD.t88 2.22001
R485 VDD.n5 VDD.t79 2.22001
R486 VDD.n64 VDD.t103 2.15435
R487 VDD.n64 VDD.t35 2.15435
R488 VDD.n37 VDD.t145 2.10455
R489 VDD.n37 VDD.t86 2.10455
R490 VDD.n36 VDD.t125 2.10455
R491 VDD.n36 VDD.t81 2.10455
R492 VDD.n2 VDD.t50 2.10455
R493 VDD.n2 VDD.t85 2.10455
R494 VDD.n3 VDD.t152 2.06607
R495 VDD.n11 VDD.t12 1.931
R496 VDD.n100 VDD.t161 1.84822
R497 VDD.n100 VDD.t45 1.84822
R498 VDD.n65 VDD.t159 1.84822
R499 VDD.n65 VDD.t37 1.84822
R500 VDD.n6 VDD.t11 1.67844
R501 VDD.n3 VDD.t150 1.4923
R502 VDD.n8 VDD.t15 1.4923
R503 VDD.n8 VDD.t3 1.4923
R504 VDD.n9 VDD.t7 1.4923
R505 VDD.n9 VDD.t17 1.4923
R506 VDD.n12 VDD.t5 1.4923
R507 VDD.n12 VDD.t13 1.4923
R508 VDD.n58 VDD.n57 1.14644
R509 VDD.n34 VDD.n33 1.14644
R510 VDD.n117 VDD.n116 1.1255
R511 VDD.n59 VDD.n34 0.9215
R512 VDD.n59 VDD.n58 0.563
R513 VDD.n97 VDD.n96 0.563
R514 VDD.n97 VDD.n59 0.359
R515 VDD.n103 VDD.n102 0.35675
R516 VDD.n117 VDD.n97 0.342875
R517 VDD.n104 VDD.n103 0.3365
R518 VDD.n102 VDD.n101 0.3065
R519 VDD.n112 VDD.n111 0.3065
R520 VDD.n110 VDD.n109 0.3065
R521 VDD.n108 VDD.n107 0.3065
R522 VDD.n50 VDD.n49 0.305021
R523 VDD.n51 VDD.n50 0.2705
R524 VDD.n107 VDD.n106 0.26
R525 VDD.n21 VDD.n20 0.149678
R526 VDD.n48 VDD.n47 0.142281
R527 VDD.n113 VDD.n104 0.1415
R528 VDD.n113 VDD.n112 0.14075
R529 VDD.n20 VDD.n19 0.131185
R530 VDD.n74 VDD.n73 0.126253
R531 VDD.n52 VDD.n51 0.120089
R532 VDD.n72 VDD.n71 0.115158
R533 VDD.n111 VDD.n110 0.1145
R534 VDD.n109 VDD.n108 0.1145
R535 VDD.n53 VDD.n52 0.113925
R536 VDD.n23 VDD.n22 0.113925
R537 VDD.n115 VDD.n99 0.109611
R538 VDD.n49 VDD.n48 0.10776
R539 VDD.n16 VDD.n15 0.106527
R540 VDD.n88 VDD.n87 0.103753
R541 VDD.n18 VDD.n17 0.100363
R542 VDD.n25 VDD.n24 0.0929658
R543 VDD.n81 VDD.n80 0.0920411
R544 VDD.n77 VDD.n76 0.080637
R545 VDD.n106 VDD.n105 0.07775
R546 VDD.n28 VDD.n27 0.0757055
R547 VDD.n27 VDD.n26 0.0744726
R548 VDD.n90 VDD.n89 0.0723151
R549 VDD.n85 VDD.n84 0.0692329
R550 VDD.n24 VDD.n23 0.0646096
R551 VDD.n54 VDD.n53 0.0624521
R552 VDD.n30 VDD.n29 0.0624521
R553 VDD.n69 VDD.n68 0.0584452
R554 VDD.n76 VDD.n75 0.0584452
R555 VDD.n78 VDD.n77 0.0584452
R556 VDD.n84 VDD.n83 0.0575205
R557 VDD.n46 VDD.n45 0.0559795
R558 VDD.n70 VDD.n69 0.0501233
R559 VDD.n83 VDD.n82 0.0473493
R560 VDD.n86 VDD.n85 0.0473493
R561 VDD.n80 VDD.n79 0.0470411
R562 VDD.n26 VDD.n25 0.0461164
R563 VDD.n57 VDD.n56 0.0456716
R564 VDD.n33 VDD.n32 0.0456716
R565 VDD.n116 VDD.n98 0.04025
R566 VDD.n17 VDD.n16 0.0387192
R567 VDD.n29 VDD.n28 0.0387192
R568 VDD.n89 VDD.n88 0.0353288
R569 VDD.n82 VDD.n81 0.0347123
R570 VDD.n94 VDD.n92 0.0331712
R571 VDD.n15 VDD.n14 0.0325548
R572 VDD.n91 VDD.n90 0.0322466
R573 VDD.n55 VDD.n54 0.0322466
R574 VDD.n31 VDD.n30 0.0322466
R575 VDD.n22 VDD.n21 0.0251575
R576 VDD.n93 VDD.n61 0.0239247
R577 VDD.n14 VDD.n13 0.0239247
R578 VDD.n87 VDD.n86 0.023
R579 VDD.n96 VDD.n60 0.0168356
R580 VDD.n96 VDD.n95 0.0168356
R581 VDD.n58 VDD.n35 0.0168356
R582 VDD.n34 VDD.n0 0.0168356
R583 VDD.n71 VDD.n70 0.0115959
R584 VDD.n73 VDD.n72 0.0115959
R585 VDD.n79 VDD.n78 0.0115959
R586 VDD VDD.n117 0.0108125
R587 VDD.n75 VDD.n74 0.0100548
R588 VDD.n19 VDD.n18 0.00789726
R589 VDD.n47 VDD.n46 0.00296575
R590 VDD.n105 VDD.n99 0.00275
R591 VDD.n92 VDD.n91 0.00142466
R592 VDD.n94 VDD.n93 0.00142466
R593 VDD.n56 VDD.n55 0.00142466
R594 VDD.n32 VDD.n31 0.00142466
R595 F6.n6 F6.n5 7.13263
R596 F6.n6 F6.n4 6.43746
R597 F6.n12 F6.n1 6.43746
R598 F6.n11 F6.n3 6.43746
R599 F6.n5 F6.t0 3.8098
R600 F6.n5 F6.t2 3.8098
R601 F6.n4 F6.t1 3.8098
R602 F6.n4 F6.t3 3.8098
R603 F6.n1 F6.t6 3.8098
R604 F6.n1 F6.t4 3.8098
R605 F6.n3 F6.t5 3.8098
R606 F6.n3 F6.t7 3.8098
R607 F6.n9 F6.n8 3.34593
R608 F6.n9 F6.n7 2.71593
R609 F6.n12 F6.n0 2.71593
R610 F6.n11 F6.n2 2.71593
R611 F6.n7 F6.t15 2.06607
R612 F6.n7 F6.t14 2.06607
R613 F6.n8 F6.t8 2.06607
R614 F6.n8 F6.t12 2.06607
R615 F6.n0 F6.t11 2.06607
R616 F6.n0 F6.t9 2.06607
R617 F6.n2 F6.t13 2.06607
R618 F6.n2 F6.t10 2.06607
R619 F6.n10 F6.n6 0.382224
R620 F6.n10 F6.n9 0.346437
R621 F6.n12 F6.n11 0.138582
R622 F6.n11 F6.n10 0.0627603
R623 F6 F6.n12 0.00173288
R624 a_484_n4228.n2 a_484_n4228.t7 121.874
R625 a_484_n4228.t7 a_484_n4228.t3 61.5152
R626 a_484_n4228.n0 a_484_n4228.t2 52.378
R627 a_484_n4228.n0 a_484_n4228.t4 17.7882
R628 a_484_n4228.n1 a_484_n4228.t0 11.1158
R629 a_484_n4228.n1 a_484_n4228.n2 9.95623
R630 a_484_n4228.n1 a_484_n4228.n0 8.37615
R631 a_484_n4228.t1 a_484_n4228.n1 8.02846
R632 a_484_n4228.n0 a_484_n4228.t6 7.3005
R633 a_484_n4228.n2 a_484_n4228.t5 6.7165
R634 a_484_n3673.n2 a_484_n3673.t6 121.874
R635 a_484_n3673.t6 a_484_n3673.t2 61.5152
R636 a_484_n3673.n0 a_484_n3673.t7 52.378
R637 a_484_n3673.n0 a_484_n3673.t5 17.7152
R638 a_484_n3673.n1 a_484_n3673.t0 11.1158
R639 a_484_n3673.n1 a_484_n3673.n2 9.95623
R640 a_484_n3673.n1 a_484_n3673.n0 8.37615
R641 a_484_n3673.t1 a_484_n3673.n1 8.02846
R642 a_484_n3673.n0 a_484_n3673.t4 7.36133
R643 a_484_n3673.n2 a_484_n3673.t3 6.7165
R644 a_757_n1888.t0 a_757_n1888.n1 21.2275
R645 a_757_n1888.n1 a_757_n1888.t4 18.9805
R646 a_757_n1888.n0 a_757_n1888.t5 17.5205
R647 a_757_n1888.n0 a_757_n1888.t2 11.5588
R648 a_757_n1888.n1 a_757_n1888.t3 11.4372
R649 a_757_n1888.t0 a_757_n1888.t1 8.60523
R650 a_757_n1888.t0 a_757_n1888.n0 8.27396
R651 VCOIN.n1 VCOIN.t2 28.7301
R652 VCOIN.n0 VCOIN.t1 18.7615
R653 VCOIN.n0 VCOIN.t0 13.5055
R654 VCOIN VCOIN.n1 5.03916
R655 VCOIN.n1 VCOIN.n0 1.01439
R656 UP UP.t0 10.0811
R657 UP UP.t1 4.27633
R658 DOWN DOWN.t0 10.0811
R659 DOWN DOWN.t1 4.27633
R660 CLK.n0 CLK.t1 17.5205
R661 CLK.n0 CLK.t0 11.5588
R662 CLK CLK.n0 11.0313
C0 a_124_n2844 a_1877_n1888 0.235746f
C1 a_673_472 a_3024_472 0.041108f
C2 a_2752_n2359 a_1332_n2408 0.014406f
C3 a_1452_n2315 a_1824_n2359 0.107446f
C4 VDD a_896_n4641 1.11099f
C5 a_1824_n3709 a_1332_n2408 0.026991f
C6 a_124_n2844 a_896_n2729 0.090966f
C7 VDD a_1804_n496 0.204841f
C8 a_1317_24 a_757_24 0.061398f
C9 VDD a_1824_n4271 0.186107f
C10 VDD a_3956_n3352 0.222895f
C11 a_2459_n3297 a_1332_n2408 0.051285f
C12 a_2576_472 a_3024_472 0.480927f
C13 a_1332_n3709 a_1332_n2408 0.154909f
C14 a_1317_n1888 a_1877_n1888 0.542819f
C15 VCOIN a_124_n4756 0.010026f
C16 VDD a_4044_n3449 0.336735f
C17 a_372_n404 a_820_n404 0.012222f
C18 VDD a_2752_n4271 0.524797f
C19 a_757_24 a_1877_n1888 0.46019f
C20 a_1356_n496 a_1268_n404 0.285629f
C21 VDD a_372_n404 0.346078f
C22 VDD a_1452_n2315 0.400846f
C23 VDD CLK 0.731835f
C24 VDD a_1233_n1440 1.07274f
C25 a_1452_n3665 a_1332_n2408 0.045667f
C26 a_224_n1440 a_673_n1440 0.051973f
C27 VDD a_673_n1440 1.4854f
C28 a_1877_n1888 a_3703_n1844 0.010209f
C29 a_673_472 a_1233_n1440 0.173051f
C30 a_2459_n2683 a_896_n2729 0.416346f
C31 a_124_n2844 a_1317_n1888 0.060492f
C32 a_224_n2800 a_896_n2729 0.071077f
C33 VDD a_1452_n4227 0.397859f
C34 a_673_472 a_673_n1440 0.01764f
C35 a_1317_24 a_1356_n496 0.010389f
C36 a_124_n2844 a_2459_n2683 0.042898f
C37 a_372_n404 a_460_n496 0.285629f
C38 a_124_n2844 a_224_n2800 0.77448f
C39 VDD a_896_n3352 1.1139f
C40 a_2752_n3709 a_1332_n2408 0.24646f
C41 a_1716_n404 a_1356_n496 0.086905f
C42 a_2576_n1440 a_1877_n1888 0.051499f
C43 VDD a_4044_n2408 0.133852f
C44 VDD a_2164_n404 0.340986f
C45 VDD a_3956_n4228 0.361712f
C46 VDD a_2459_n4595 0.371422f
C47 VDD a_2752_n2359 0.523241f
C48 a_1877_n1888 a_3024_n1440 0.057075f
C49 VDD a_1824_n3709 0.186132f
C50 a_896_n2729 a_1332_n2408 0.280621f
C51 a_n76_n404 a_372_n404 0.012222f
C52 VDD a_1233_472 0.996523f
C53 a_1332_n3709 a_1792_n5184 0.016718f
C54 VDD a_2459_n3297 0.370377f
C55 a_124_n2844 a_1332_n2408 0.137044f
C56 VDD a_1332_n3709 0.58464f
C57 a_1268_n404 a_820_n404 0.012552f
C58 a_1824_n4271 a_896_n4641 1.16391f
C59 VDD a_3956_n2316 0.355683f
C60 VDD a_224_472 0.460056f
C61 a_673_472 a_1233_472 0.79492f
C62 VDD a_1268_n404 0.336412f
C63 a_673_472 a_224_472 0.051973f
C64 a_36_n3352 a_36_n4712 0.010569f
C65 VDD a_1452_n3665 0.397896f
C66 a_896_n4641 a_2752_n4271 0.023074f
C67 VDD a_36_n3352 0.278953f
C68 VDD a_1317_24 0.472916f
C69 a_896_n2729 a_1824_n2359 1.16391f
C70 a_3956_n3352 a_4044_n3449 0.285629f
C71 a_908_n496 a_1268_n404 0.086905f
C72 VDD a_1716_n404 0.332254f
C73 VDD a_12_n496 0.254868f
C74 a_2576_472 a_1233_472 0.097396f
C75 a_124_n2844 a_1824_n2359 0.032377f
C76 VDD a_2752_n3709 0.520925f
C77 a_1317_24 a_673_472 0.318865f
C78 a_224_n5184 VCOIN 0.455456f
C79 a_2459_n2683 a_1332_n2408 0.011266f
C80 a_1792_n5184 F6 1.62795f
C81 a_1452_n4227 a_896_n4641 0.839895f
C82 VDD F6 0.818211f
C83 a_224_n2800 a_1332_n2408 0.107397f
C84 VDD a_1877_n1888 1.78852f
C85 a_1824_n4271 a_1452_n4227 0.107446f
C86 a_896_n4641 a_2459_n4595 0.416346f
C87 a_12_n496 a_460_n496 0.013276f
C88 a_673_472 a_1877_n1888 0.290117f
C89 a_2164_n404 a_1804_n496 0.086905f
C90 VDD a_896_n2729 1.11698f
C91 VDD a_124_n3449 0.377703f
C92 a_3024_472 a_1233_472 0.224841f
C93 a_2576_n1440 a_3024_n1440 0.480927f
C94 a_673_n1440 a_1233_n1440 0.77678f
C95 a_224_n1440 a_124_n2844 0.517726f
C96 a_1824_n4271 a_2459_n4595 0.021118f
C97 a_36_n4712 a_124_n4756 0.285629f
C98 VDD a_124_n2844 1.49699f
C99 a_2459_n2683 a_1824_n2359 0.021118f
C100 VDD VCOIN 0.658453f
C101 VDD a_124_n4756 0.377188f
C102 a_1332_n3709 a_896_n4641 0.093423f
C103 a_2576_472 a_1877_n1888 0.050704f
C104 a_2752_n4271 a_2459_n4595 0.493186f
C105 a_n76_n404 a_12_n496 0.285629f
C106 DOWN a_1877_n1888 0.01269f
C107 a_2164_n404 a_673_n1440 0.019418f
C108 a_1332_n3709 a_1824_n4271 0.046461f
C109 VDD a_1317_n1888 0.472672f
C110 VDD a_2459_n2683 0.372354f
C111 VDD a_757_24 1.81567f
C112 VDD a_224_n2800 0.827537f
C113 a_1332_n2408 a_1824_n2359 0.018863f
C114 a_1332_n3709 a_2752_n4271 0.266557f
C115 a_3956_n2316 a_4044_n3449 0.010569f
C116 a_1233_472 a_1233_n1440 0.013905f
C117 a_3024_472 a_1877_n1888 0.05477f
C118 a_673_472 a_757_24 0.776323f
C119 CLK a_224_472 0.502436f
C120 a_1716_n404 a_1804_n496 0.285629f
C121 a_896_n3352 a_1824_n3709 1.16391f
C122 VDD a_2252_n496 0.231745f
C123 VDD a_4044_n4320 0.131342f
C124 a_1332_n3709 a_1452_n4227 0.032472f
C125 UP a_757_24 0.473919f
C126 VDD a_2576_n1440 0.57564f
C127 a_1877_n1888 a_1804_n496 0.014853f
C128 a_896_n3352 a_2459_n3297 0.416346f
C129 a_896_n3352 a_1332_n3709 0.307596f
C130 a_2576_472 a_757_24 0.036901f
C131 a_1332_n3709 a_3956_n4228 0.025816f
C132 VDD a_1332_n2408 1.21408f
C133 a_4044_n2408 a_3956_n2316 0.285629f
C134 VDD a_3024_n1440 0.443621f
C135 a_372_n404 a_12_n496 0.086742f
C136 a_2752_n3709 a_2752_n4271 0.01024f
C137 a_1332_n3709 a_2459_n4595 0.05056f
C138 VDD a_1356_n496 0.208364f
C139 a_2459_n3297 a_1824_n3709 0.021118f
C140 a_1716_n404 a_673_n1440 0.011215f
C141 a_896_n3352 a_1452_n3665 0.839895f
C142 a_1332_n3709 a_1824_n3709 0.01975f
C143 a_1877_n1888 a_3703_68 0.010314f
C144 a_1877_n1888 a_1233_n1440 0.870988f
C145 a_1877_n1888 a_673_n1440 0.131931f
C146 a_896_n3352 a_2752_n3709 0.023074f
C147 a_1332_n3709 a_2459_n3297 0.010957f
C148 a_908_n496 a_1356_n496 0.013276f
C149 a_1824_n3709 a_1452_n3665 0.107446f
C150 a_2164_n404 a_1716_n404 0.012552f
C151 a_896_n2729 a_1452_n2315 0.839895f
C152 a_3024_472 a_757_24 0.048924f
C153 VDD a_224_n5184 1.01168f
C154 VDD a_1824_n2359 0.186856f
C155 a_124_n2844 a_1452_n2315 0.025834f
C156 a_673_n1440 a_896_n2729 0.010446f
C157 a_896_n4641 a_224_n2800 0.421686f
C158 a_1332_n3709 a_1452_n3665 0.242122f
C159 a_124_n2844 a_673_n1440 0.029378f
C160 a_1317_24 a_1233_472 0.827579f
C161 a_2459_n3297 a_2752_n3709 0.493186f
C162 a_1332_n3709 a_2752_n3709 0.015243f
C163 a_1716_n404 a_1268_n404 0.012552f
C164 VDD a_36_n4712 0.278953f
C165 a_896_n2729 a_2752_n2359 0.023074f
C166 a_1804_n496 a_2252_n496 0.013276f
C167 VDD a_820_n404 0.343186f
C168 VDD a_1792_n5184 1.90337f
C169 VDD a_224_n1440 0.465743f
C170 a_1317_n1888 a_1233_n1440 0.827579f
C171 a_1233_472 a_1877_n1888 1.28745f
C172 a_124_n2844 a_2752_n2359 0.249206f
C173 a_1317_n1888 a_673_n1440 0.318976f
C174 VDD a_673_472 1.25124f
C175 CLK a_757_24 0.020177f
C176 a_4044_n4320 a_3956_n3352 0.010569f
C177 a_820_n404 a_460_n496 0.086742f
C178 a_908_n496 a_820_n404 0.285629f
C179 VDD a_460_n496 0.215083f
C180 VDD UP 0.129208f
C181 a_1356_n496 a_1804_n496 0.013276f
C182 VDD a_908_n496 0.211978f
C183 a_3956_n3352 a_1332_n2408 0.023971f
C184 a_1452_n4227 a_224_n2800 0.227561f
C185 a_3956_n2316 a_124_n2844 0.026006f
C186 a_2252_n496 a_673_n1440 0.026153f
C187 a_1317_24 a_1877_n1888 0.542819f
C188 a_896_n3352 a_224_n2800 0.075252f
C189 a_2576_n1440 a_1233_n1440 0.099075f
C190 VDD a_2576_472 0.565435f
C191 a_4044_n3449 a_1332_n2408 0.010299f
C192 VDD DOWN 0.129208f
C193 a_36_n3352 a_124_n3449 0.285629f
C194 a_2459_n2683 a_2752_n2359 0.493186f
C195 a_2576_n1440 a_673_n1440 0.524f
C196 a_1452_n2315 a_1332_n2408 0.240887f
C197 a_2576_472 a_673_472 0.524441f
C198 a_908_n496 a_460_n496 0.013276f
C199 a_3024_n1440 a_1233_n1440 0.232395f
C200 a_2164_n404 a_2252_n496 0.285629f
C201 VDD a_n76_n404 0.404801f
C202 a_4044_n4320 a_3956_n4228 0.285629f
C203 a_1233_472 a_757_24 0.590855f
C204 VDD a_3024_472 0.436971f
C205 a_896_n3352 a_1332_n2408 0.098711f
C206 a_1332_n3709 a_224_n2800 0.147928f
C207 a_224_472 a_757_24 0.259946f
C208 F6 GND 1.07141f
C209 VCOIN GND 0.726876f
C210 DOWN GND 0.219834f
C211 UP GND 0.190568f
C212 CLK GND 0.578798f
C213 VDD GND 57.681072f
C214 a_1792_n5184 GND 3.00173f
C215 a_224_n5184 GND 1.55349f
C216 a_3956_n4228 GND 0.356232f
C217 a_4044_n4320 GND 0.615444f
C218 a_2459_n4595 GND 0.469002f
C219 a_2752_n4271 GND 0.85819f
C220 a_1452_n4227 GND 0.304138f
C221 a_1824_n4271 GND 0.42522f
C222 a_896_n4641 GND 1.48203f
C223 a_124_n4756 GND 0.253352f
C224 a_36_n4712 GND 0.509546f
C225 a_3956_n3352 GND 0.555186f
C226 a_4044_n3449 GND 0.3597f
C227 a_2752_n3709 GND 0.858306f
C228 a_2459_n3297 GND 0.469151f
C229 a_1452_n3665 GND 0.304138f
C230 a_1824_n3709 GND 0.42522f
C231 a_1332_n3709 GND 1.37227f
C232 a_896_n3352 GND 1.48111f
C233 a_36_n3352 GND 0.509546f
C234 a_124_n3449 GND 0.255426f
C235 a_3956_n2316 GND 0.355739f
C236 a_4044_n2408 GND 0.623811f
C237 a_2459_n2683 GND 0.474447f
C238 a_2752_n2359 GND 0.862377f
C239 a_1452_n2315 GND 0.30791f
C240 a_1824_n2359 GND 0.425059f
C241 a_1332_n2408 GND 0.699352f
C242 a_896_n2729 GND 1.48407f
C243 a_224_n2800 GND 0.744772f
C244 a_3024_n1440 GND 0.504963f
C245 a_2576_n1440 GND 0.529868f
C246 a_1317_n1888 GND 0.653228f
C247 a_224_n1440 GND 0.48757f
C248 a_124_n2844 GND 2.4228f
C249 a_1233_n1440 GND 1.35363f
C250 a_673_n1440 GND 1.62629f
C251 a_2164_n404 GND 0.291705f
C252 a_1716_n404 GND 0.285378f
C253 a_1268_n404 GND 0.286621f
C254 a_820_n404 GND 0.288647f
C255 a_372_n404 GND 0.288752f
C256 a_n76_n404 GND 0.290611f
C257 a_2252_n496 GND 0.497887f
C258 a_1804_n496 GND 0.476784f
C259 a_1356_n496 GND 0.479397f
C260 a_908_n496 GND 0.484202f
C261 a_460_n496 GND 0.483304f
C262 a_12_n496 GND 0.494234f
C263 a_3024_472 GND 0.510031f
C264 a_2576_472 GND 0.536139f
C265 a_1877_n1888 GND 3.92094f
C266 a_1233_472 GND 1.42826f
C267 a_1317_24 GND 0.668914f
C268 a_673_472 GND 1.94746f
C269 a_757_24 GND 1.54832f
C270 a_224_472 GND 0.496642f
C271 a_757_n1888.t0 GND 1.25053f
C272 a_757_n1888.t1 GND 0.048467f
C273 a_757_n1888.t5 GND 0.077986f
C274 a_757_n1888.t2 GND 0.042413f
C275 a_757_n1888.n0 GND 0.079885f
C276 a_757_n1888.t4 GND 0.078379f
C277 a_757_n1888.t3 GND 0.060967f
C278 a_757_n1888.n1 GND 0.46137f
C279 a_484_n3673.t4 GND 0.042682f
C280 a_484_n3673.n0 GND 0.221505f
C281 a_484_n3673.n1 GND 0.803219f
C282 a_484_n3673.t2 GND 0.127787f
C283 a_484_n3673.t6 GND 0.401653f
C284 a_484_n3673.t3 GND 0.020325f
C285 a_484_n3673.n2 GND 0.257957f
C286 a_484_n3673.t7 GND 0.144509f
C287 a_484_n3673.t5 GND 0.127878f
C288 a_484_n3673.t0 GND 0.047684f
C289 a_484_n3673.t1 GND 0.1048f
C290 a_484_n4228.t6 GND 0.043151f
C291 a_484_n4228.n0 GND 0.221428f
C292 a_484_n4228.n1 GND 0.803219f
C293 a_484_n4228.t2 GND 0.144509f
C294 a_484_n4228.t4 GND 0.127487f
C295 a_484_n4228.t0 GND 0.047684f
C296 a_484_n4228.t5 GND 0.020325f
C297 a_484_n4228.t3 GND 0.127787f
C298 a_484_n4228.t7 GND 0.401653f
C299 a_484_n4228.n2 GND 0.257957f
C300 a_484_n4228.t1 GND 0.1048f
C301 VDD.n0 GND 0.025629f
C302 VDD.t139 GND 0.074279f
C303 VDD.t8 GND 0.156005f
C304 VDD.t111 GND 0.052431f
C305 VDD.t4 GND 0.070911f
C306 VDD.t12 GND 0.044266f
C307 VDD.t155 GND 0.032373f
C308 VDD.t141 GND 0.048134f
C309 VDD.t143 GND 0.089821f
C310 VDD.t84 GND 0.055869f
C311 VDD.t147 GND 0.043836f
C312 VDD.t49 GND 0.048134f
C313 VDD.t149 GND 0.055869f
C314 VDD.t151 GND 0.085094f
C315 VDD.t137 GND 0.048134f
C316 VDD.t153 GND 0.030728f
C317 VDD.n10 GND 0.107491f
C318 VDD.t76 GND 0.015901f
C319 VDD.t99 GND 0.032662f
C320 VDD.t165 GND 0.051572f
C321 VDD.t78 GND 0.046415f
C322 VDD.t126 GND 0.043836f
C323 VDD.t87 GND 0.06425f
C324 VDD.t108 GND 0.052431f
C325 VDD.t82 GND 0.056944f
C326 VDD.t10 GND 0.055869f
C327 VDD.t136 GND 0.037819f
C328 VDD.t134 GND 0.048134f
C329 VDD.t2 GND 0.053291f
C330 VDD.t28 GND 0.043836f
C331 VDD.t14 GND 0.057589f
C332 VDD.t16 GND 0.069622f
C333 VDD.t132 GND 0.043836f
C334 VDD.t6 GND 0.078647f
C335 VDD.n11 GND 0.057837f
C336 VDD.n13 GND 0.074267f
C337 VDD.n14 GND 0.013036f
C338 VDD.n15 GND 0.041115f
C339 VDD.n16 GND 0.030479f
C340 VDD.n17 GND 0.032939f
C341 VDD.n18 GND 0.023211f
C342 VDD.n19 GND 0.030768f
C343 VDD.n20 GND 0.056464f
C344 VDD.n21 GND 0.036293f
C345 VDD.n22 GND 0.032209f
C346 VDD.n23 GND 0.037609f
C347 VDD.n24 GND 0.036241f
C348 VDD.n25 GND 0.03225f
C349 VDD.n26 GND 0.025633f
C350 VDD.n27 GND 0.033142f
C351 VDD.n28 GND 0.024018f
C352 VDD.n29 GND 0.025959f
C353 VDD.n30 GND 0.018644f
C354 VDD.n33 GND 0.209774f
C355 VDD.n34 GND 0.117139f
C356 VDD.n35 GND 0.025629f
C357 VDD.t30 GND 0.074279f
C358 VDD.t109 GND 0.100565f
C359 VDD.t80 GND 0.133657f
C360 VDD.t124 GND 0.136665f
C361 VDD.t121 GND 0.123558f
C362 VDD.t63 GND 0.067046f
C363 VDD.n42 GND 0.082248f
C364 VDD.t48 GND 0.047704f
C365 VDD.t24 GND 0.078217f
C366 VDD.t20 GND 0.110665f
C367 VDD.t123 GND 0.125492f
C368 VDD.t120 GND 0.094763f
C369 VDD.t68 GND 0.086813f
C370 VDD.t89 GND 0.12807f
C371 VDD.t70 GND 0.151707f
C372 VDD.n43 GND 0.084052f
C373 VDD.t46 GND 0.252702f
C374 VDD.n44 GND 0.078466f
C375 VDD.n45 GND 0.081575f
C376 VDD.n46 GND 0.025368f
C377 VDD.n47 GND 0.042327f
C378 VDD.n48 GND 0.060549f
C379 VDD.n49 GND 0.088184f
C380 VDD.n50 GND 0.123045f
C381 VDD.n51 GND 0.086789f
C382 VDD.n52 GND 0.053444f
C383 VDD.n53 GND 0.040737f
C384 VDD.n54 GND 0.018644f
C385 VDD.n55 GND 0.012728f
C386 VDD.n57 GND 0.209774f
C387 VDD.n58 GND 0.031725f
C388 VDD.n59 GND 0.514732f
C389 VDD.n60 GND 0.025629f
C390 VDD.n61 GND 0.166955f
C391 VDD.t61 GND 0.064992f
C392 VDD.t32 GND 0.096268f
C393 VDD.t115 GND 0.096482f
C394 VDD.t128 GND 0.057374f
C395 VDD.t97 GND 0.08273f
C396 VDD.t59 GND 0.076498f
C397 VDD.t91 GND 0.081441f
C398 VDD.t18 GND 0.058663f
C399 VDD.t53 GND 0.076498f
C400 VDD.t38 GND 0.096268f
C401 VDD.t51 GND 0.043836f
C402 VDD.t162 GND 0.071341f
C403 VDD.n62 GND 0.092433f
C404 VDD.t117 GND 0.062316f
C405 VDD.t93 GND 0.071341f
C406 VDD.n63 GND 0.101673f
C407 VDD.t106 GND 0.068977f
C408 VDD.t95 GND 0.050498f
C409 VDD.t34 GND 0.087672f
C410 VDD.t102 GND 0.051572f
C411 VDD.t22 GND 0.043836f
C412 VDD.t42 GND 0.043836f
C413 VDD.t36 GND 0.051572f
C414 VDD.t158 GND 0.056514f
C415 VDD.n66 GND 0.066602f
C416 VDD.t72 GND 0.051712f
C417 VDD.n67 GND 0.068042f
C418 VDD.n68 GND 0.213089f
C419 VDD.n69 GND 0.035119f
C420 VDD.n70 GND 0.014664f
C421 VDD.n71 GND 0.027629f
C422 VDD.n72 GND 0.030705f
C423 VDD.n73 GND 0.028547f
C424 VDD.n74 GND 0.029506f
C425 VDD.n75 GND 0.019571f
C426 VDD.n76 GND 0.041115f
C427 VDD.n77 GND 0.033441f
C428 VDD.n78 GND 0.027549f
C429 VDD.n79 GND 0.017601f
C430 VDD.n80 GND 0.033225f
C431 VDD.n81 GND 0.030986f
C432 VDD.n82 GND 0.022021f
C433 VDD.n83 GND 0.026503f
C434 VDD.n84 GND 0.030986f
C435 VDD.n85 GND 0.028804f
C436 VDD.n86 GND 0.019719f
C437 VDD.n87 GND 0.030986f
C438 VDD.n88 GND 0.033225f
C439 VDD.n89 GND 0.027231f
C440 VDD.n90 GND 0.020582f
C441 VDD.n91 GND 0.012728f
C442 VDD.n93 GND 0.01106f
C443 VDD.n95 GND 0.025671f
C444 VDD.n97 GND 0.372154f
C445 VDD.n98 GND 0.010512f
C446 VDD.t55 GND 0.114855f
C447 VDD.t160 GND 0.059415f
C448 VDD.t44 GND 0.043836f
C449 VDD.t0 GND 0.072953f
C450 VDD.t65 GND 0.099168f
C451 VDD.t100 GND 0.079292f
C452 VDD.n101 GND 0.053378f
C453 VDD.n102 GND 0.027972f
C454 VDD.n103 GND 0.029281f
C455 VDD.n104 GND 0.022138f
C456 VDD.n106 GND 0.011291f
C457 VDD.n107 GND 0.024859f
C458 VDD.n108 GND 0.02003f
C459 VDD.n109 GND 0.02003f
C460 VDD.n110 GND 0.02003f
C461 VDD.n111 GND 0.02003f
C462 VDD.n112 GND 0.020901f
C463 VDD.n113 GND 0.023316f
C464 VDD.n114 GND 0.067614f
C465 VDD.t156 GND 0.052969f
C466 VDD.t40 GND 0.060167f
C467 VDD.t113 GND 0.060167f
C468 VDD.t104 GND 0.060167f
C469 VDD.t57 GND 0.060167f
C470 VDD.t26 GND 0.070159f
C471 VDD.t130 GND 0.080009f
C472 VDD.n115 GND 0.102597f
C473 VDD.n116 GND 0.01299f
C474 VDD.n117 GND 0.187272f
C475 a_484_n2316.t2 GND 0.041275f
C476 a_484_n2316.n0 GND 0.211801f
C477 a_484_n2316.n1 GND 0.768297f
C478 a_484_n2316.t4 GND 0.138226f
C479 a_484_n2316.t5 GND 0.121944f
C480 a_484_n2316.t0 GND 0.045611f
C481 a_484_n2316.t7 GND 0.019441f
C482 a_484_n2316.t6 GND 0.122231f
C483 a_484_n2316.t3 GND 0.38419f
C484 a_484_n2316.n2 GND 0.246741f
C485 a_484_n2316.t1 GND 0.100244f
C486 a_572_n4284.n0 GND 0.686004f
C487 a_572_n4284.t3 GND 0.024037f
C488 a_572_n4284.t2 GND 0.019883f
C489 a_572_n4284.n1 GND 1.27029f
C490 a_572_n4284.t0 GND 0.067797f
C491 a_572_n4284.t1 GND 0.063309f
C492 a_572_n4284.t11 GND 0.052652f
C493 a_572_n4284.t6 GND 0.034715f
C494 a_572_n4284.t7 GND 0.019483f
C495 a_572_n4284.n2 GND 0.092881f
C496 a_572_n4284.t16 GND 0.034715f
C497 a_572_n4284.t4 GND 0.019483f
C498 a_572_n4284.n3 GND 0.060005f
C499 a_572_n4284.t15 GND 0.034715f
C500 a_572_n4284.t8 GND 0.019483f
C501 a_572_n4284.t13 GND 0.024223f
C502 a_572_n4284.t14 GND 0.025812f
C503 a_572_n4284.n4 GND 0.056612f
C504 a_572_n4284.t10 GND 0.025916f
C505 a_572_n4284.t5 GND 0.024113f
C506 a_572_n4284.n5 GND 0.046919f
C507 a_572_n4284.t9 GND 0.024223f
C508 a_572_n4284.t12 GND 0.025812f
C509 a_572_n4284.n6 GND 0.046914f
.ends

