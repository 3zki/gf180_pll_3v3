* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt cp_layout CSVB UP DOWN VCNB VCNS OUT GND VDD
X0 VDD.t34 a_373_1386.t3 a_2144_800 VDD.t33 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X1 a_3208_800 a_373_1386.t4 VDD.t32 VDD.t31 pfet_03v3 ad=0.52p pd=2.52u as=1.3p ps=5.3u w=2u l=0.33u
X2 a_543_1260.t0 VCNB.t4 a_3944_0 GND.t37 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X3 OUT.t7 a_1398_660 a_614_800 VDD.t24 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X4 OUT.t1 DOWN.t0 a_614_0 GND.t1 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X5 a_444_800 a_373_1386.t5 VDD.t30 VDD.t29 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X6 VDD.t2 UP.t0 a_1398_660 VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0.52p ps=2.52u w=2u l=0.33u
X7 a_3208_800 a_543_1260.t3 a_373_1386.t0 VDD.t13 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X8 OUT.t3 DOWN.t1 a_614_0 GND.t11 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X9 GND.t9 VCNS.t4 a_3208_0 GND.t8 nfet_03v3 ad=0.4p pd=1.8u as=0.26p ps=1.52u w=1u l=0.33u
X10 a_373_1386.t0 a_543_1260.t4 a_3208_800 VDD.t15 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X11 VDD.t12 CSVB.t0 VCNB.t0 VDD.t11 pfet_03v3 ad=1.456p pd=5.78u as=0.5824p ps=2.76u w=2.24u l=0.56u
X12 VDD.t26 DOWN.t2 a_104_0 VDD.t25 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X13 a_614_800 a_1398_660 OUT.t6 VDD.t23 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X14 a_1398_660 UP.t1 VDD.t10 VDD.t9 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X15 a_614_0 VCNB.t5 a_444_0 GND.t36 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X16 a_614_0 a_104_0 a_784_0 GND.t27 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X17 VDD.t28 a_373_1386.t6 a_3208_800 VDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.52p ps=2.52u w=2u l=0.33u
X18 GND.t21 UP.t2 a_1398_660 GND.t20 nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.33u
X19 a_614_800 a_543_1260.t5 a_444_800 VDD.t0 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X20 a_543_1260.t2 a_543_1260.t1 VDD.t20 VDD.t19 pfet_03v3 ad=1.072p pd=5.3u as=1.072p ps=5.3u w=0.8u l=0.33u
X21 a_3208_0 VCNS.t5 GND.t17 GND.t16 nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.33u
X22 GND.t23 VCNS.t6 a_5008_0 GND.t22 nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.33u
X23 VCNB.t3 VCNB.t2 GND.t35 GND.t34 nfet_03v3 ad=0.496p pd=3.22u as=0.496p ps=3.22u w=0.4u l=0.33u
X24 a_614_800 UP.t3 a_784_0 VDD.t5 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X25 a_1398_660 UP.t4 GND.t41 GND.t40 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X26 a_104_0 DOWN.t3 VDD.t4 VDD.t3 pfet_03v3 ad=0.52p pd=2.52u as=1.3p ps=5.3u w=2u l=0.33u
X27 a_2144_0 VCNB.t6 a_614_0 GND.t33 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X28 GND.t5 VCNS.t7 a_3944_0 GND.t4 nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.33u
X29 a_784_0 UP.t5 a_614_800 VDD.t8 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X30 a_3944_0 VCNB.t7 a_543_1260.t0 GND.t32 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X31 a_5008_0 VCNS.t8 GND.t13 GND.t12 nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.33u
X32 a_614_0 DOWN.t4 OUT.t0 GND.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X33 VCNS.t3 CSVB.t1 VDD.t37 VDD.t36 pfet_03v3 ad=0.5824p pd=2.76u as=1.456p ps=5.78u w=2.24u l=0.56u
X34 a_3944_0 VCNS.t9 GND.t7 GND.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.4p ps=1.8u w=1u l=0.33u
X35 a_784_0 UP.t6 a_614_800 VDD.t14 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X36 a_614_0 a_104_0 a_784_0 GND.t26 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X37 a_614_0 DOWN.t5 OUT.t2 GND.t10 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X38 a_784_0 a_104_0 a_614_0 GND.t25 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X39 OUT.t5 a_1398_660 a_614_800 VDD.t22 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X40 VCNB.t1 CSVB.t2 VDD.t17 VDD.t16 pfet_03v3 ad=0.5824p pd=2.76u as=0.5824p ps=2.76u w=2.24u l=0.56u
X41 a_3208_0 VCNB.t8 a_373_1386.t1 GND.t31 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X42 a_444_0 VCNS.t10 GND.t15 GND.t14 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X43 a_784_0 a_104_0 a_614_0 GND.t24 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X44 VDD.t7 CSVB.t3 VCNS.t0 VDD.t6 pfet_03v3 ad=0.5824p pd=2.76u as=0.5824p ps=2.76u w=2.24u l=0.56u
X45 a_373_1386.t2 VCNB.t9 a_3208_0 GND.t30 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X46 a_614_800 UP.t7 a_784_0 VDD.t18 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X47 a_104_0 DOWN.t6 GND.t39 GND.t38 nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.33u
X48 GND.t19 DOWN.t7 a_104_0 GND.t18 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X49 a_5008_0 VCNB.t10 VCNS.t2 GND.t29 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X50 a_614_800 a_1398_660 OUT.t4 VDD.t21 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X51 a_2144_800 a_543_1260.t6 a_614_800 VDD.t35 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X52 GND.t3 VCNS.t11 a_2144_0 GND.t2 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
X53 VCNS.t1 VCNB.t11 a_5008_0 GND.t28 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.33u
R0 a_373_1386.n0 a_373_1386.t5 56.5589
R1 a_373_1386.n1 a_373_1386.t6 54.6191
R2 a_373_1386.n1 a_373_1386.t4 54.3444
R3 a_373_1386.n0 a_373_1386.t3 54.3444
R4 a_373_1386.n3 a_373_1386.n2 7.32981
R5 a_373_1386.n3 a_373_1386.n1 3.5139
R6 a_373_1386.t0 a_373_1386.n3 1.76266
R7 a_373_1386.n2 a_373_1386.t1 1.6385
R8 a_373_1386.n2 a_373_1386.t2 1.6385
R9 a_373_1386.n1 a_373_1386.n0 1.33205
R10 VDD.n3 VDD.t11 494.065
R11 VDD.n8 VDD.t36 480.769
R12 VDD.n18 VDD.t3 457.205
R13 VDD.t19 VDD.n8 443.911
R14 VDD.n9 VDD.t19 443.911
R15 VDD.n9 VDD.t27 443.911
R16 VDD.n17 VDD.t31 443.911
R17 VDD.t1 VDD.n17 443.911
R18 VDD.t11 VDD.t16 346.154
R19 VDD.t16 VDD.t6 346.154
R20 VDD.t6 VDD.t36 346.154
R21 VDD.t27 VDD.t13 272.437
R22 VDD.t13 VDD.t15 272.437
R23 VDD.t15 VDD.t31 272.437
R24 VDD.t9 VDD.t1 272.437
R25 VDD.t33 VDD.t9 272.437
R26 VDD.t35 VDD.t33 272.437
R27 VDD.t23 VDD.t35 272.437
R28 VDD.t24 VDD.t23 272.437
R29 VDD.t21 VDD.t24 272.437
R30 VDD.t22 VDD.t21 272.437
R31 VDD.t18 VDD.t22 272.437
R32 VDD.t14 VDD.t18 272.437
R33 VDD.t5 VDD.t14 272.437
R34 VDD.t8 VDD.t5 272.437
R35 VDD.t0 VDD.t8 272.437
R36 VDD.t29 VDD.t0 272.437
R37 VDD.t25 VDD.t29 272.437
R38 VDD.t3 VDD.t25 272.437
R39 VDD.n2 VDD.t20 14.4695
R40 VDD.n17 VDD.n16 13.2611
R41 VDD.n10 VDD.n9 13.2611
R42 VDD.n8 VDD.n7 13.2611
R43 VDD.n18 VDD.t4 12.2645
R44 VDD.n15 VDD.t2 12.2645
R45 VDD.n12 VDD.t32 12.2645
R46 VDD.n11 VDD.t28 12.2645
R47 VDD.n1 VDD.n0 10.7945
R48 VDD.n14 VDD.n13 10.7945
R49 VDD.n6 VDD.t37 9.44208
R50 VDD.n3 VDD.t12 9.44208
R51 VDD.n5 VDD.n4 8.12958
R52 VDD.n0 VDD.t30 0.9105
R53 VDD.n0 VDD.t26 0.9105
R54 VDD.n13 VDD.t10 0.9105
R55 VDD.n13 VDD.t34 0.9105
R56 VDD.n4 VDD.t17 0.813
R57 VDD.n4 VDD.t7 0.813
R58 VDD.n14 VDD.n1 0.437643
R59 VDD.n12 VDD.n11 0.159929
R60 VDD.n5 VDD.n3 0.0999286
R61 VDD.n6 VDD.n5 0.0999286
R62 VDD.n7 VDD.n2 0.0849286
R63 VDD.n15 VDD.n14 0.0802143
R64 VDD VDD.n1 0.0617857
R65 VDD.n7 VDD.n6 0.0347857
R66 VDD.n10 VDD.n2 0.0347857
R67 VDD.n11 VDD.n10 0.0347857
R68 VDD.n16 VDD.n12 0.0347857
R69 VDD.n16 VDD.n15 0.0347857
R70 VDD VDD.n18 0.0189286
R71 VCNB.n10 VCNB.t5 29.3475
R72 VCNB.n9 VCNB.t6 29.3475
R73 VCNB.n8 VCNB.t9 29.3475
R74 VCNB.n7 VCNB.t8 29.3475
R75 VCNB.n6 VCNB.t4 29.3475
R76 VCNB.n5 VCNB.t7 29.3475
R77 VCNB.n4 VCNB.t11 29.3475
R78 VCNB.n3 VCNB.t10 29.3475
R79 VCNB.n2 VCNB.t2 29.3475
R80 VCNB.n1 VCNB.t3 10.616
R81 VCNB.n1 VCNB.n0 2.94063
R82 VCNB.n10 VCNB.n9 1.81234
R83 VCNB.n9 VCNB.n8 1.46182
R84 VCNB.n5 VCNB.n4 1.05918
R85 VCNB.n0 VCNB.t0 0.813
R86 VCNB.n0 VCNB.t1 0.813
R87 VCNB VCNB.n10 0.778526
R88 VCNB.n7 VCNB.n6 0.670763
R89 VCNB.n3 VCNB.n2 0.649447
R90 VCNB.n2 VCNB.n1 0.321421
R91 VCNB.n4 VCNB.n3 0.201816
R92 VCNB.n6 VCNB.n5 0.201816
R93 VCNB.n8 VCNB.n7 0.201816
R94 a_543_1260.n0 a_543_1260.t5 42.2199
R95 a_543_1260.n0 a_543_1260.t6 40.4081
R96 a_543_1260.n0 a_543_1260.t4 40.4081
R97 a_543_1260.n0 a_543_1260.t3 40.4081
R98 a_543_1260.n1 a_543_1260.t1 40.4081
R99 a_543_1260.t0 a_543_1260.n1 7.4853
R100 a_543_1260.n1 a_543_1260.t2 5.40883
R101 a_543_1260.n1 a_543_1260.n0 2.96695
R102 GND.t22 GND.t34 1323.81
R103 GND.t34 GND.n4 994.173
R104 GND.n16 GND.t38 994.072
R105 GND.n5 GND.t12 970.097
R106 GND.n5 GND.t4 970.097
R107 GND.n15 GND.t16 970.097
R108 GND.t20 GND.n15 970.097
R109 GND.t6 GND.t8 791.487
R110 GND.t29 GND.t22 595.366
R111 GND.t28 GND.t29 595.366
R112 GND.t12 GND.t28 595.366
R113 GND.t4 GND.t32 595.366
R114 GND.t32 GND.t37 595.366
R115 GND.t37 GND.t6 595.366
R116 GND.t8 GND.t31 595.366
R117 GND.t31 GND.t30 595.366
R118 GND.t30 GND.t16 595.366
R119 GND.t40 GND.t20 595.366
R120 GND.t2 GND.t40 595.366
R121 GND.t33 GND.t2 595.366
R122 GND.t0 GND.t33 595.366
R123 GND.t1 GND.t0 595.366
R124 GND.t10 GND.t1 595.366
R125 GND.t11 GND.t10 595.366
R126 GND.t27 GND.t11 595.366
R127 GND.t24 GND.t27 595.366
R128 GND.t26 GND.t24 595.366
R129 GND.t25 GND.t26 595.366
R130 GND.t36 GND.t25 595.366
R131 GND.t14 GND.t36 595.366
R132 GND.t18 GND.t14 595.366
R133 GND.t38 GND.t18 595.366
R134 GND.n4 GND.t35 24.116
R135 GND.n6 GND.n5 23.9005
R136 GND.n15 GND.n14 23.9005
R137 GND.n16 GND.t39 22.3205
R138 GND.n13 GND.t21 22.3205
R139 GND.n10 GND.t17 22.3205
R140 GND.n7 GND.t5 22.3205
R141 GND.n2 GND.t13 22.3205
R142 GND.n3 GND.t23 22.3205
R143 GND.n1 GND.n0 19.8005
R144 GND.n12 GND.n11 19.8005
R145 GND.n9 GND.n8 19.8005
R146 GND.n8 GND.t7 2.5205
R147 GND.n8 GND.t9 2.5205
R148 GND.n0 GND.t15 1.6385
R149 GND.n0 GND.t19 1.6385
R150 GND.n11 GND.t41 1.6385
R151 GND.n11 GND.t3 1.6385
R152 GND.n12 GND.n1 0.9185
R153 GND.n3 GND.n2 0.3317
R154 GND.n9 GND.n7 0.3317
R155 GND.n10 GND.n9 0.3317
R156 GND.n13 GND.n12 0.1661
R157 GND GND.n16 0.0887
R158 GND GND.n1 0.0779
R159 GND.n6 GND.n2 0.0743
R160 GND.n7 GND.n6 0.0743
R161 GND.n14 GND.n10 0.0743
R162 GND.n14 GND.n13 0.0743
R163 GND.n4 GND.n3 0.0689
R164 OUT.n3 OUT.n2 11.4305
R165 OUT OUT.n5 11.1943
R166 OUT.n4 OUT.n0 4.27695
R167 OUT.n3 OUT.n1 4.27695
R168 OUT.n5 OUT.t0 1.6385
R169 OUT.n5 OUT.t1 1.6385
R170 OUT.n2 OUT.t2 1.6385
R171 OUT.n2 OUT.t3 1.6385
R172 OUT.n0 OUT.t6 0.9105
R173 OUT.n0 OUT.t7 0.9105
R174 OUT.n1 OUT.t4 0.9105
R175 OUT.n1 OUT.t5 0.9105
R176 OUT.n4 OUT.n3 0.383
R177 OUT OUT.n4 0.23675
R178 DOWN.n3 DOWN.t2 47.5611
R179 DOWN.n4 DOWN.t7 36.5005
R180 DOWN.n1 DOWN.t1 33.21
R181 DOWN.n0 DOWN.t4 33.21
R182 DOWN.n3 DOWN.t3 28.7581
R183 DOWN.n5 DOWN.n3 26.2141
R184 DOWN.n4 DOWN.t6 17.6975
R185 DOWN.n1 DOWN.t5 17.6975
R186 DOWN.n0 DOWN.t0 17.6975
R187 DOWN.n5 DOWN.n4 10.7293
R188 DOWN.n6 DOWN.n5 8.0005
R189 DOWN.n2 DOWN.n0 7.75675
R190 DOWN.n2 DOWN.n1 7.75675
R191 DOWN.n6 DOWN.n2 3.21483
R192 DOWN DOWN.n6 0.04325
R193 UP.n3 UP.t1 47.5611
R194 UP.n0 UP.t7 44.2706
R195 UP.n1 UP.t5 44.2706
R196 UP.n4 UP.t4 36.5005
R197 UP.n3 UP.t0 28.7581
R198 UP.n0 UP.t6 28.7581
R199 UP.n1 UP.t3 28.7581
R200 UP.n5 UP.n4 26.2141
R201 UP.n4 UP.t2 17.6975
R202 UP.n5 UP.n3 10.7293
R203 UP.n6 UP.n5 9.54625
R204 UP.n2 UP.n0 7.75675
R205 UP.n2 UP.n1 7.75675
R206 UP.n6 UP.n2 1.66908
R207 UP UP.n6 1.382
R208 VCNS.n3 VCNS.t6 43.5585
R209 VCNS.n10 VCNS.t10 43.2838
R210 VCNS.n9 VCNS.t11 43.2838
R211 VCNS.n8 VCNS.t5 43.2838
R212 VCNS.n7 VCNS.t4 43.2838
R213 VCNS.n6 VCNS.t9 43.2838
R214 VCNS.n5 VCNS.t7 43.2838
R215 VCNS.n4 VCNS.t8 43.2838
R216 VCNS.n2 VCNS.n1 6.3005
R217 VCNS.n3 VCNS.n2 5.67959
R218 VCNS.n2 VCNS.n0 2.56843
R219 VCNS.n10 VCNS.n9 2.21497
R220 VCNS.n1 VCNS.t2 1.6385
R221 VCNS.n1 VCNS.t1 1.6385
R222 VCNS.n9 VCNS.n8 1.05918
R223 VCNS.n0 VCNS.t0 0.813
R224 VCNS.n0 VCNS.t3 0.813
R225 VCNS.n5 VCNS.n4 0.654303
R226 VCNS.n6 VCNS.n5 0.604447
R227 VCNS.n8 VCNS.n7 0.604447
R228 VCNS VCNS.n10 0.577211
R229 VCNS.n4 VCNS.n3 0.275613
R230 VCNS.n7 VCNS.n6 0.268132
R231 CSVB.n0 CSVB.t1 29.2438
R232 CSVB CSVB.t0 29.1266
R233 CSVB.n0 CSVB.t3 28.988
R234 CSVB.n1 CSVB.t2 28.988
R235 CSVB.n1 CSVB.n0 0.256289
R236 CSVB CSVB.n1 0.117737
C0 a_5008_0 VCNB 0.210175f
C1 VDD VCNB 0.469741f
C2 DOWN UP 1.44253f
C3 DOWN VCNB 0.146186f
C4 VCNS a_5008_0 0.510902f
C5 a_614_800 OUT 1.18823f
C6 VCNS VDD 0.381004f
C7 VDD OUT 0.036564f
C8 VCNS DOWN 0.021642f
C9 DOWN OUT 0.209353f
C10 a_3208_800 VDD 0.702282f
C11 a_614_800 a_614_0 0.145142f
C12 a_104_0 a_784_0 0.24687f
C13 CSVB VCNB 0.149254f
C14 DOWN a_614_0 0.110426f
C15 a_2144_800 a_1398_660 0.012025f
C16 a_5008_0 VDD 0.018357f
C17 VCNS CSVB 0.158612f
C18 a_614_800 VDD 0.580264f
C19 a_1398_660 UP 1.42689f
C20 a_104_0 UP 0.091313f
C21 a_784_0 UP 0.32679f
C22 a_614_800 DOWN 0.016002f
C23 DOWN VDD 0.306675f
C24 VCNB a_1398_660 0.038456f
C25 a_3944_0 VCNB 0.200645f
C26 a_104_0 VCNB 0.203456f
C27 VCNB a_784_0 0.076741f
C28 OUT a_1398_660 0.305455f
C29 VCNS a_3944_0 0.038289f
C30 VCNS a_104_0 0.018945f
C31 a_784_0 OUT 0.109016f
C32 VCNB UP 0.063044f
C33 VCNB a_3208_0 0.200558f
C34 VCNS UP 0.022937f
C35 OUT UP 0.112163f
C36 VCNS VCNB 6.34632f
C37 VCNB OUT 0.075053f
C38 VCNS a_3208_0 0.038289f
C39 a_5008_0 CSVB 0.014166f
C40 CSVB VDD 0.738439f
C41 a_104_0 a_614_0 0.111757f
C42 a_784_0 a_614_0 0.394051f
C43 a_614_800 a_1398_660 0.186658f
C44 VDD a_1398_660 1.06596f
C45 a_3944_0 VDD 0.036853f
C46 a_614_800 a_784_0 1.15373f
C47 a_104_0 VDD 0.512285f
C48 VDD a_784_0 0.039903f
C49 a_614_0 UP 0.031663f
C50 a_614_800 a_2144_800 0.019086f
C51 VDD a_2144_800 0.02646f
C52 DOWN a_1398_660 0.023562f
C53 a_3208_800 a_3208_0 0.062097f
C54 VCNB a_614_0 0.223159f
C55 a_104_0 DOWN 1.41006f
C56 DOWN a_784_0 0.10389f
C57 a_614_800 a_444_800 0.019086f
C58 VDD a_444_800 0.02646f
C59 VCNS a_614_0 0.033577f
C60 OUT a_614_0 0.36483f
C61 a_614_800 UP 0.211047f
C62 VDD UP 0.869486f
C63 VCNB GND 3.950222f
C64 VCNS GND 4.249971f
C65 OUT GND 0.203842f
C66 CSVB GND 0.759737f
C67 UP GND 1.51484f
C68 DOWN GND 1.86882f
C69 VDD GND 14.1656f
C70 a_5008_0 GND 0.69875f
C71 a_3944_0 GND 0.714938f
C72 a_3208_0 GND 0.695632f
C73 a_2144_0 GND 0.012152f
C74 a_614_0 GND 0.735429f
C75 a_444_0 GND 0.012152f
C76 a_3208_800 GND 0.092226f
C77 a_784_0 GND 0.18513f
C78 a_614_800 GND 0.286671f
C79 a_104_0 GND 1.23694f
C80 a_1398_660 GND 0.673787f
C81 VCNS.t0 GND 0.081375f
C82 VCNS.t3 GND 0.081375f
C83 VCNS.n0 GND 0.366808f
C84 VCNS.t2 GND 0.036328f
C85 VCNS.t1 GND 0.036328f
C86 VCNS.n1 GND 0.072657f
C87 VCNS.n2 GND 0.686508f
C88 VCNS.t6 GND 0.110829f
C89 VCNS.n3 GND 0.737889f
C90 VCNS.t8 GND 0.109584f
C91 VCNS.n4 GND 0.324673f
C92 VCNS.t7 GND 0.109584f
C93 VCNS.n5 GND 0.358978f
C94 VCNS.t9 GND 0.109584f
C95 VCNS.n6 GND 0.272338f
C96 VCNS.t4 GND 0.109584f
C97 VCNS.n7 GND 0.272338f
C98 VCNS.t5 GND 0.109584f
C99 VCNS.n8 GND 0.449676f
C100 VCNS.t11 GND 0.109584f
C101 VCNS.n9 GND 0.810724f
C102 VCNS.t10 GND 0.109584f
C103 VCNS.n10 GND 0.702675f
C104 a_543_1260.t0 GND 0.197147f
C105 a_543_1260.n0 GND 2.37979f
C106 a_543_1260.n1 GND 1.01023f
C107 a_543_1260.t5 GND 0.187773f
C108 a_543_1260.t6 GND 0.151828f
C109 a_543_1260.t4 GND 0.151828f
C110 a_543_1260.t3 GND 0.151828f
C111 a_543_1260.t1 GND 0.040321f
C112 a_543_1260.t2 GND 0.029257f
C113 VCNB.t0 GND 0.088433f
C114 VCNB.t1 GND 0.088433f
C115 VCNB.n0 GND 0.486426f
C116 VCNB.t3 GND 0.099496f
C117 VCNB.n1 GND 0.821119f
C118 VCNB.t2 GND 0.027866f
C119 VCNB.n2 GND 0.300642f
C120 VCNB.t10 GND 0.087995f
C121 VCNB.n3 GND 0.25872f
C122 VCNB.t11 GND 0.087995f
C123 VCNB.n4 GND 0.358541f
C124 VCNB.t7 GND 0.087995f
C125 VCNB.n5 GND 0.358541f
C126 VCNB.t4 GND 0.087995f
C127 VCNB.n6 GND 0.263913f
C128 VCNB.t8 GND 0.087995f
C129 VCNB.n7 GND 0.263913f
C130 VCNB.t9 GND 0.087995f
C131 VCNB.n8 GND 0.45663f
C132 VCNB.t6 GND 0.087995f
C133 VCNB.n9 GND 0.848989f
C134 VCNB.t5 GND 0.087995f
C135 VCNB.n10 GND 0.682525f
C136 a_373_1386.t0 GND 0.261348f
C137 a_373_1386.n0 GND 1.48854f
C138 a_373_1386.n1 GND 1.07597f
C139 a_373_1386.t1 GND 0.032497f
C140 a_373_1386.t2 GND 0.032497f
C141 a_373_1386.n2 GND 0.096598f
C142 a_373_1386.t6 GND 0.161342f
C143 a_373_1386.t5 GND 0.190482f
C144 a_373_1386.t3 GND 0.160334f
C145 a_373_1386.t4 GND 0.160334f
C146 a_373_1386.n3 GND 0.640059f
.ends

